library verilog;
use verilog.vl_types.all;
entity stoplight is
    port(
        reset_n         : in     vl_logic;
        clk             : in     vl_logic;
        northsouth_red  : out    vl_logic;
        northsouth_yellow: out    vl_logic;
        northsouth_green: out    vl_logic;
        eastwest_red    : out    vl_logic;
        eastwest_yellow : out    vl_logic;
        eastwest_green  : out    vl_logic
    );
end stoplight;
