
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, n6, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ns;

  DFFARX1 \reg_b_reg[0]  ( .D(N92), .CLK(clk), .RSTB(n331), .Q(reg_b[0]), .QN(
        n252) );
  DFFARX1 \reg_a_reg[4]  ( .D(N63), .CLK(clk), .RSTB(n328), .QN(n217) );
  DFFARX1 \reg_b_reg[5]  ( .D(N97), .CLK(clk), .RSTB(n329), .Q(n106), .QN(n220) );
  DFFARX1 \reg_b_reg[1]  ( .D(N93), .CLK(clk), .RSTB(n331), .Q(reg_b[1]), .QN(
        n223) );
  DFFARX1 \reg_a_reg[6]  ( .D(N65), .CLK(clk), .RSTB(n329), .QN(n140) );
  DFFARX1 \reg_a_reg[5]  ( .D(N64), .CLK(clk), .RSTB(n329), .QN(n139) );
  DFFARX1 \gcd_ps_reg[0]  ( .D(gcd_ns[0]), .CLK(clk), .RSTB(n332), .Q(n191), 
        .QN(n67) );
  DFFARX1 \reg_a_reg[20]  ( .D(N79), .CLK(clk), .RSTB(n322), .Q(reg_a[20]), 
        .QN(n161) );
  DFFARX1 \gcd_ps_reg[1]  ( .D(gcd_ns[1]), .CLK(clk), .RSTB(n331), .Q(n209), 
        .QN(n100) );
  DFFARX1 \reg_a_reg[13]  ( .D(N72), .CLK(clk), .RSTB(n318), .Q(reg_a[13]), 
        .QN(n165) );
  DFFARX1 \reg_b_reg[29]  ( .D(N121), .CLK(clk), .RSTB(n326), .Q(reg_b[29]), 
        .QN(n201) );
  DFFARX1 \reg_b_reg[30]  ( .D(N122), .CLK(clk), .RSTB(n327), .Q(reg_b[30]), 
        .QN(n202) );
  DFFARX1 \reg_a_reg[3]  ( .D(N62), .CLK(clk), .RSTB(n328), .Q(reg_a[3]), .QN(
        n164) );
  DFFARX1 \reg_a_reg[19]  ( .D(N78), .CLK(clk), .RSTB(n321), .Q(reg_a[19]), 
        .QN(n159) );
  DFFARX1 \reg_a_reg[16]  ( .D(N75), .CLK(clk), .RSTB(n320), .Q(reg_a[16]), 
        .QN(n166) );
  DFFARX1 \reg_a_reg[21]  ( .D(N80), .CLK(clk), .RSTB(n322), .Q(reg_a[21]), 
        .QN(n200) );
  DFFARX1 \reg_a_reg[12]  ( .D(N71), .CLK(clk), .RSTB(n318), .Q(reg_a[12]), 
        .QN(n203) );
  DFFARX1 \reg_a_reg[18]  ( .D(N77), .CLK(clk), .RSTB(n321), .Q(reg_a[18]), 
        .QN(n198) );
  DFFARX1 \reg_a_reg[24]  ( .D(N83), .CLK(clk), .RSTB(n324), .Q(reg_a[24]), 
        .QN(n197) );
  DFFARX1 \reg_a_reg[15]  ( .D(N74), .CLK(clk), .RSTB(n319), .Q(reg_a[15]), 
        .QN(n199) );
  DFFARX1 \reg_b_reg[25]  ( .D(N117), .CLK(clk), .RSTB(n324), .Q(reg_b[25]), 
        .QN(n205) );
  DFFARX1 \reg_b_reg[21]  ( .D(N113), .CLK(clk), .RSTB(n322), .Q(reg_b[21]), 
        .QN(n206) );
  DFFARX1 \reg_b_reg[10]  ( .D(N102), .CLK(clk), .RSTB(n317), .Q(reg_b[10]), 
        .QN(n204) );
  DFFARX1 \reg_b_reg[18]  ( .D(N110), .CLK(clk), .RSTB(n321), .Q(reg_b[18]), 
        .QN(n193) );
  DFFARX1 \reg_b_reg[22]  ( .D(N114), .CLK(clk), .RSTB(n323), .Q(reg_b[22]), 
        .QN(n208) );
  DFFARX1 \reg_b_reg[24]  ( .D(N116), .CLK(clk), .RSTB(n324), .Q(reg_b[24]), 
        .QN(n196) );
  DFFARX1 \reg_b_reg[19]  ( .D(N111), .CLK(clk), .RSTB(n321), .Q(reg_b[19]), 
        .QN(n195) );
  DFFARX1 \reg_b_reg[15]  ( .D(N107), .CLK(clk), .RSTB(n319), .Q(reg_b[15]), 
        .QN(n192) );
  DFFARX1 \reg_b_reg[16]  ( .D(N108), .CLK(clk), .RSTB(n320), .Q(reg_b[16]), 
        .QN(n157) );
  DFFARX1 \reg_b_reg[9]  ( .D(N101), .CLK(clk), .RSTB(n316), .Q(reg_b[9]), 
        .QN(n207) );
  DFFARX1 \reg_b_reg[12]  ( .D(N104), .CLK(clk), .RSTB(n318), .Q(reg_b[12]), 
        .QN(n194) );
  DFFARX1 \reg_a_reg[28]  ( .D(N87), .CLK(clk), .RSTB(n326), .Q(reg_a[28]), 
        .QN(n190) );
  DFFARX1 \reg_a_reg[31]  ( .D(N90), .CLK(clk), .RSTB(n330), .Q(reg_a[31]), 
        .QN(n155) );
  DFFARX1 \reg_b_reg[2]  ( .D(N94), .CLK(clk), .RSTB(n327), .Q(reg_b[2]), .QN(
        n189) );
  DFFARX1 \reg_b_reg[8]  ( .D(N100), .CLK(clk), .RSTB(n316), .Q(reg_b[8]), 
        .QN(n125) );
  DFFARX1 \reg_a_reg[1]  ( .D(N60), .CLK(clk), .RSTB(n331), .QN(n146) );
  DFFARX1 \reg_b_reg[6]  ( .D(N98), .CLK(clk), .RSTB(n329), .Q(n116), .QN(n215) );
  DFFARX1 \result_reg[31]  ( .D(n97), .CLK(clk), .RSTB(n330), .Q(result[31])
         );
  DFFARX1 \result_reg[7]  ( .D(n96), .CLK(clk), .RSTB(n330), .Q(result[7]) );
  DFFARX1 \result_reg[1]  ( .D(n98), .CLK(clk), .RSTB(n331), .Q(result[1]) );
  DFFARX1 \result_reg[8]  ( .D(n68), .CLK(clk), .RSTB(n316), .Q(result[8]) );
  DFFARX1 \result_reg[20]  ( .D(n80), .CLK(clk), .RSTB(n322), .Q(result[20])
         );
  DFFARX1 \result_reg[19]  ( .D(n79), .CLK(clk), .RSTB(n321), .Q(result[19])
         );
  DFFARX1 \result_reg[18]  ( .D(n78), .CLK(clk), .RSTB(n321), .Q(result[18])
         );
  DFFARX1 \result_reg[17]  ( .D(n77), .CLK(clk), .RSTB(n320), .Q(result[17])
         );
  DFFARX1 \result_reg[16]  ( .D(n76), .CLK(clk), .RSTB(n320), .Q(result[16])
         );
  DFFARX1 \result_reg[15]  ( .D(n75), .CLK(clk), .RSTB(n319), .Q(result[15])
         );
  DFFARX1 \result_reg[14]  ( .D(n74), .CLK(clk), .RSTB(n319), .Q(result[14])
         );
  DFFARX1 \result_reg[13]  ( .D(n73), .CLK(clk), .RSTB(n318), .Q(result[13])
         );
  DFFARX1 \result_reg[12]  ( .D(n72), .CLK(clk), .RSTB(n318), .Q(result[12])
         );
  DFFARX1 \result_reg[11]  ( .D(n71), .CLK(clk), .RSTB(n317), .Q(result[11])
         );
  DFFARX1 \result_reg[10]  ( .D(n70), .CLK(clk), .RSTB(n317), .Q(result[10])
         );
  DFFARX1 \result_reg[9]  ( .D(n69), .CLK(clk), .RSTB(n316), .Q(result[9]) );
  DFFARX1 \result_reg[30]  ( .D(n90), .CLK(clk), .RSTB(n327), .Q(result[30])
         );
  DFFARX1 \result_reg[29]  ( .D(n89), .CLK(clk), .RSTB(n326), .Q(result[29])
         );
  DFFARX1 \result_reg[28]  ( .D(n88), .CLK(clk), .RSTB(n326), .Q(result[28])
         );
  DFFARX1 \result_reg[27]  ( .D(n87), .CLK(clk), .RSTB(n325), .Q(result[27])
         );
  DFFARX1 \result_reg[26]  ( .D(n86), .CLK(clk), .RSTB(n325), .Q(result[26])
         );
  DFFARX1 \result_reg[25]  ( .D(n85), .CLK(clk), .RSTB(n324), .Q(result[25])
         );
  DFFARX1 \result_reg[24]  ( .D(n84), .CLK(clk), .RSTB(n324), .Q(result[24])
         );
  DFFARX1 \result_reg[23]  ( .D(n83), .CLK(clk), .RSTB(n323), .Q(result[23])
         );
  DFFARX1 \result_reg[22]  ( .D(n82), .CLK(clk), .RSTB(n323), .Q(result[22])
         );
  DFFARX1 \result_reg[21]  ( .D(n81), .CLK(clk), .RSTB(n322), .Q(result[21])
         );
  DFFARX1 \result_reg[6]  ( .D(n95), .CLK(clk), .RSTB(n329), .Q(result[6]) );
  DFFARX1 \result_reg[5]  ( .D(n94), .CLK(clk), .RSTB(n329), .Q(result[5]) );
  DFFARX1 \result_reg[4]  ( .D(n93), .CLK(clk), .RSTB(n328), .Q(result[4]) );
  DFFARX1 \result_reg[3]  ( .D(n92), .CLK(clk), .RSTB(n328), .Q(result[3]) );
  DFFARX1 \result_reg[2]  ( .D(n91), .CLK(clk), .RSTB(n327), .Q(result[2]) );
  DFFARX1 \result_reg[0]  ( .D(n99), .CLK(clk), .RSTB(n331), .Q(result[0]) );
  DFFARX1 \reg_a_reg[26]  ( .D(N85), .CLK(clk), .RSTB(n325), .Q(reg_a[26]), 
        .QN(n511) );
  DFFARX1 \reg_b_reg[4]  ( .D(N96), .CLK(clk), .RSTB(n328), .Q(n105), .QN(n218) );
  DFFARX1 \reg_b_reg[28]  ( .D(N120), .CLK(clk), .RSTB(n326), .Q(reg_b[28]) );
  DFFARX1 \reg_b_reg[31]  ( .D(N123), .CLK(clk), .RSTB(n330), .Q(reg_b[31]), 
        .QN(n563) );
  DFFARX1 \reg_b_reg[20]  ( .D(N112), .CLK(clk), .RSTB(n322), .Q(reg_b[20]), 
        .QN(n346) );
  DFFARX1 \reg_b_reg[27]  ( .D(N119), .CLK(clk), .RSTB(n325), .Q(reg_b[27]) );
  DFFARX1 \reg_b_reg[13]  ( .D(N105), .CLK(clk), .RSTB(n318), .Q(reg_b[13]), 
        .QN(n355) );
  DFFARX1 \reg_b_reg[26]  ( .D(N118), .CLK(clk), .RSTB(n325), .Q(reg_b[26]), 
        .QN(n342) );
  DFFARX1 \reg_b_reg[23]  ( .D(N115), .CLK(clk), .RSTB(n323), .Q(reg_b[23]), 
        .QN(n343) );
  DFFARX1 \reg_b_reg[17]  ( .D(N109), .CLK(clk), .RSTB(n320), .Q(reg_b[17]), 
        .QN(n349) );
  DFFARX1 \reg_b_reg[14]  ( .D(N106), .CLK(clk), .RSTB(n319), .Q(reg_b[14]), 
        .QN(n352) );
  DFFARX1 \reg_b_reg[11]  ( .D(N103), .CLK(clk), .RSTB(n317), .Q(reg_b[11]), 
        .QN(n356) );
  DFFARX1 \reg_b_reg[3]  ( .D(N95), .CLK(clk), .RSTB(n328), .Q(reg_b[3]) );
  DFFARX1 \reg_a_reg[22]  ( .D(N81), .CLK(clk), .RSTB(n323), .Q(reg_a[22]) );
  DFFARX1 \reg_a_reg[23]  ( .D(N82), .CLK(clk), .RSTB(n323), .Q(reg_a[23]) );
  DFFARX1 \reg_a_reg[27]  ( .D(N86), .CLK(clk), .RSTB(n325), .Q(reg_a[27]), 
        .QN(n398) );
  DFFARX1 \reg_a_reg[11]  ( .D(N70), .CLK(clk), .RSTB(n317), .Q(reg_a[11]) );
  DFFARX1 \reg_a_reg[10]  ( .D(N69), .CLK(clk), .RSTB(n317), .Q(reg_a[10]) );
  DFFARX1 \reg_a_reg[17]  ( .D(N76), .CLK(clk), .RSTB(n320), .Q(reg_a[17]) );
  DFFARX1 \reg_a_reg[14]  ( .D(N73), .CLK(clk), .RSTB(n319), .Q(reg_a[14]) );
  DFFARX1 \reg_a_reg[30]  ( .D(N89), .CLK(clk), .RSTB(n327), .Q(reg_a[30]) );
  DFFARX1 \reg_a_reg[29]  ( .D(N88), .CLK(clk), .RSTB(n326), .Q(reg_a[29]) );
  DFFARX1 \reg_a_reg[25]  ( .D(N84), .CLK(clk), .RSTB(n324), .Q(reg_a[25]) );
  DFFARX1 \reg_a_reg[9]  ( .D(N68), .CLK(clk), .RSTB(n316), .Q(reg_a[9]) );
  DFFARX1 \reg_a_reg[8]  ( .D(N67), .CLK(clk), .RSTB(n316), .Q(reg_a[8]) );
  DFFARX1 \reg_a_reg[7]  ( .D(N66), .CLK(clk), .RSTB(n330), .Q(reg_a[7]) );
  DFFARX1 \reg_b_reg[7]  ( .D(N99), .CLK(clk), .RSTB(n330), .Q(reg_b[7]), .QN(
        n188) );
  DFFARX1 \reg_a_reg[2]  ( .D(N61), .CLK(clk), .RSTB(n327), .Q(reg_a[2]), .QN(
        n187) );
  DFFARX1 \reg_a_reg[0]  ( .D(N59), .CLK(clk), .RSTB(n332), .Q(reg_a[0]), .QN(
        n224) );
  INVX8 U166 ( .IN(n129), .QN(n102) );
  INVX8 U167 ( .IN(n129), .QN(n170) );
  INVX4 U168 ( .IN(n421), .QN(n103) );
  INVX8 U169 ( .IN(n103), .QN(n104) );
  INVX4 U170 ( .IN(n179), .QN(n585) );
  OR2X2 U171 ( .IN1(n576), .IN2(n413), .Q(n179) );
  OR2X1 U172 ( .IN1(reg_a[17]), .IN2(n349), .Q(n351) );
  OR2X1 U173 ( .IN1(reg_a[11]), .IN2(n356), .Q(n358) );
  OR2X1 U174 ( .IN1(n211), .IN2(n220), .Q(n370) );
  NAND2X0 U175 ( .IN1(n197), .IN2(reg_b[24]), .QN(n495) );
  INVX0 U176 ( .IN(n486), .QN(n344) );
  NAND2X0 U177 ( .IN1(n199), .IN2(reg_b[15]), .QN(n455) );
  INVX4 U178 ( .IN(n567), .QN(n581) );
  NAND2X0 U179 ( .IN1(n506), .IN2(n505), .QN(n507) );
  NAND2X1 U180 ( .IN1(n254), .IN2(n171), .QN(n219) );
  INVX2 U181 ( .IN(n536), .QN(n361) );
  OR2X1 U182 ( .IN1(reg_a[14]), .IN2(n352), .Q(n354) );
  INVX0 U183 ( .IN(n370), .QN(n359) );
  OR2X1 U184 ( .IN1(n190), .IN2(reg_b[28]), .Q(n401) );
  OR2X1 U185 ( .IN1(n368), .IN2(n419), .Q(n424) );
  INVX2 U186 ( .IN(n424), .QN(n373) );
  NOR2X0 U187 ( .IN1(n502), .IN2(n107), .QN(n390) );
  NAND2X0 U188 ( .IN1(n200), .IN2(reg_b[21]), .QN(n481) );
  OR2X1 U189 ( .IN1(reg_a[20]), .IN2(n346), .Q(n348) );
  AO22X1 U190 ( .IN1(n347), .IN2(n348), .IN3(reg_a[20]), .IN4(n346), .Q(n478)
         );
  INVX0 U191 ( .IN(n473), .QN(n347) );
  NBUFFX2 U192 ( .IN(n178), .Q(n147) );
  INVX0 U193 ( .IN(n460), .QN(n350) );
  INVX0 U194 ( .IN(n351), .QN(n384) );
  NAND2X0 U195 ( .IN1(n203), .IN2(reg_b[12]), .QN(n441) );
  INVX0 U196 ( .IN(n358), .QN(n380) );
  NAND2X0 U197 ( .IN1(n198), .IN2(reg_b[18]), .QN(n468) );
  INVX0 U198 ( .IN(n547), .QN(n371) );
  OR2X1 U199 ( .IN1(n576), .IN2(n413), .Q(n411) );
  OAI21X1 U200 ( .IN1(reg_a[7]), .IN2(n188), .IN3(n554), .QN(n419) );
  NAND2X1 U201 ( .IN1(n188), .IN2(reg_a[7]), .QN(n418) );
  NAND2X0 U202 ( .IN1(n204), .IN2(reg_a[10]), .QN(n432) );
  NOR4X0 U203 ( .IN1(n65), .IN2(n66), .IN3(n63), .IN4(n64), .QN(n167) );
  NOR4X0 U204 ( .IN1(n61), .IN2(n62), .IN3(n59), .IN4(n60), .QN(n168) );
  OA21X1 U205 ( .IN1(n110), .IN2(n531), .IN3(n530), .Q(n174) );
  INVX0 U206 ( .IN(n389), .QN(n492) );
  NAND2X0 U207 ( .IN1(n192), .IN2(reg_a[15]), .QN(n456) );
  NAND2X0 U208 ( .IN1(n193), .IN2(reg_a[18]), .QN(n469) );
  NAND2X1 U209 ( .IN1(n189), .IN2(reg_a[2]), .QN(n540) );
  AND2X1 U210 ( .IN1(n536), .IN2(n537), .Q(n180) );
  NAND2X0 U211 ( .IN1(n194), .IN2(reg_a[12]), .QN(n442) );
  NAND2X0 U212 ( .IN1(n195), .IN2(reg_a[19]), .QN(n473) );
  OAI21X1 U213 ( .IN1(reg_a[19]), .IN2(n195), .IN3(n468), .QN(n474) );
  INVX0 U214 ( .IN(n386), .QN(n475) );
  NAND2X0 U215 ( .IN1(n218), .IN2(n221), .QN(n547) );
  NOR2X0 U216 ( .IN1(n221), .IN2(n218), .QN(n153) );
  INVX2 U217 ( .IN(n139), .QN(n211) );
  INVX2 U218 ( .IN(n217), .QN(n221) );
  NAND2X2 U219 ( .IN1(n229), .IN2(n118), .QN(n129) );
  XOR3X1 U220 ( .IN1(reg_a[2]), .IN2(reg_b[2]), .IN3(n180), .Q(n538) );
  NBUFFX2 U221 ( .IN(n581), .Q(n258) );
  XOR3X1 U222 ( .IN1(reg_b[27]), .IN2(reg_a[27]), .IN3(n516), .Q(n518) );
  NAND2X0 U223 ( .IN1(n515), .IN2(n514), .QN(N85) );
  NOR2X0 U224 ( .IN1(n513), .IN2(n512), .QN(n514) );
  NAND2X0 U225 ( .IN1(n575), .IN2(n574), .QN(N60) );
  NOR2X0 U226 ( .IN1(n573), .IN2(n572), .QN(n574) );
  AND2X1 U227 ( .IN1(n186), .IN2(n576), .Q(gcd_ns[1]) );
  INVX0 U228 ( .IN(n229), .QN(n248) );
  NOR2X0 U229 ( .IN1(reg_a[26]), .IN2(n342), .QN(n107) );
  OR2X1 U230 ( .IN1(reg_b[27]), .IN2(n398), .Q(n108) );
  AOI22X1 U231 ( .IN1(n377), .IN2(n376), .IN3(reg_a[8]), .IN4(n125), .QN(n109)
         );
  INVX2 U232 ( .IN(n118), .QN(n255) );
  INVX2 U233 ( .IN(n118), .QN(n256) );
  INVX2 U234 ( .IN(n140), .QN(n216) );
  AND2X1 U235 ( .IN1(n401), .IN2(n400), .Q(n110) );
  OR2X1 U236 ( .IN1(n448), .IN2(n382), .Q(n111) );
  AND2X1 U237 ( .IN1(n251), .IN2(n348), .Q(n112) );
  AND2X1 U238 ( .IN1(n175), .IN2(n345), .Q(n113) );
  OR2X1 U239 ( .IN1(n461), .IN2(n384), .Q(n114) );
  AND2X1 U240 ( .IN1(n226), .IN2(n482), .Q(n115) );
  AND2X1 U241 ( .IN1(n132), .IN2(n496), .Q(n117) );
  NAND2X0 U242 ( .IN1(n167), .IN2(n168), .QN(n6) );
  OA21X2 U243 ( .IN1(n413), .IN2(n410), .IN3(n412), .Q(n118) );
  OR2X1 U244 ( .IN1(n438), .IN2(n381), .Q(n119) );
  OR2X1 U245 ( .IN1(n452), .IN2(n383), .Q(n120) );
  OR2X1 U246 ( .IN1(n433), .IN2(n380), .Q(n121) );
  AND2X1 U247 ( .IN1(n397), .IN2(n108), .Q(n122) );
  NBUFFX2 U248 ( .IN(n367), .Q(n124) );
  AOI22X1 U249 ( .IN1(n142), .IN2(reg_b[2]), .IN3(n579), .IN4(reg_a[2]), .QN(
        n123) );
  INVX2 U250 ( .IN(n146), .QN(n222) );
  NAND2X4 U251 ( .IN1(n389), .IN2(n117), .QN(n504) );
  INVX0 U252 ( .IN(n491), .QN(n132) );
  NAND2X4 U253 ( .IN1(n390), .IN2(n504), .QN(n391) );
  INVX2 U254 ( .IN(n118), .QN(n254) );
  NOR2X4 U255 ( .IN1(n104), .IN2(n214), .QN(n142) );
  NBUFFX2 U256 ( .IN(n567), .Q(n126) );
  INVX4 U257 ( .IN(n142), .QN(n127) );
  INVX8 U258 ( .IN(n127), .QN(n128) );
  NOR2X4 U259 ( .IN1(n118), .IN2(n104), .QN(n131) );
  OAI21X2 U260 ( .IN1(n413), .IN2(n410), .IN3(n412), .QN(n214) );
  INVX8 U261 ( .IN(n568), .QN(n130) );
  INVX8 U262 ( .IN(n568), .QN(n583) );
  NAND2X4 U263 ( .IN1(n373), .IN2(n417), .QN(n374) );
  NOR2X4 U264 ( .IN1(n178), .IN2(n136), .QN(n133) );
  NOR2X4 U265 ( .IN1(n133), .IN2(n134), .QN(n386) );
  AND2X1 U266 ( .IN1(n135), .IN2(n114), .Q(n134) );
  INVX0 U267 ( .IN(n143), .QN(n135) );
  OR2X1 U268 ( .IN1(n120), .IN2(n143), .Q(n136) );
  NAND2X0 U269 ( .IN1(n130), .IN2(n538), .QN(n137) );
  NAND2X0 U270 ( .IN1(a_in[2]), .IN2(n258), .QN(n138) );
  NAND3X0 U271 ( .IN1(n137), .IN2(n138), .IN3(n123), .QN(N61) );
  NOR2X0 U272 ( .IN1(n151), .IN2(n114), .QN(n150) );
  NOR2X0 U273 ( .IN1(n147), .IN2(n120), .QN(n151) );
  NOR2X4 U274 ( .IN1(n576), .IN2(n413), .QN(n228) );
  XOR3X2 U275 ( .IN1(n222), .IN2(n577), .IN3(reg_b[1]), .Q(n569) );
  OR2X2 U276 ( .IN1(n576), .IN2(n413), .Q(n229) );
  INVX4 U277 ( .IN(n410), .QN(n576) );
  OAI21X2 U278 ( .IN1(n222), .IN2(n223), .IN3(n577), .QN(n536) );
  NAND2X4 U279 ( .IN1(n366), .IN2(n365), .QN(n415) );
  OR2X2 U280 ( .IN1(n372), .IN2(n551), .Q(n417) );
  NAND2X4 U281 ( .IN1(n176), .IN2(n113), .QN(n389) );
  NAND2X2 U282 ( .IN1(n104), .IN2(n118), .QN(n567) );
  OR2X2 U283 ( .IN1(n216), .IN2(n215), .Q(n554) );
  NAND2X4 U284 ( .IN1(n364), .IN2(n539), .QN(n366) );
  NOR2X4 U285 ( .IN1(n363), .IN2(n362), .QN(n364) );
  NAND2X4 U286 ( .IN1(n374), .IN2(n375), .QN(n379) );
  INVX8 U287 ( .IN(n131), .QN(n141) );
  NAND2X4 U288 ( .IN1(n254), .IN2(n104), .QN(n568) );
  NOR2X4 U289 ( .IN1(n361), .IN2(n360), .QN(n363) );
  OR2X1 U290 ( .IN1(n465), .IN2(n385), .Q(n143) );
  OR2X1 U291 ( .IN1(n186), .IN2(n414), .Q(n144) );
  NOR2X4 U292 ( .IN1(n228), .IN2(n144), .QN(n421) );
  NOR2X0 U293 ( .IN1(n6), .IN2(n413), .QN(n186) );
  NAND2X4 U294 ( .IN1(n369), .IN2(n373), .QN(n375) );
  NOR2X4 U295 ( .IN1(n416), .IN2(n367), .QN(n369) );
  INVX4 U296 ( .IN(n415), .QN(n367) );
  NAND2X4 U297 ( .IN1(n397), .IN2(n108), .QN(n145) );
  NAND2X4 U298 ( .IN1(n227), .IN2(n115), .QN(n176) );
  NAND2X4 U299 ( .IN1(n386), .IN2(n112), .QN(n227) );
  INVX0 U300 ( .IN(n474), .QN(n251) );
  INVX0 U301 ( .IN(n478), .QN(n226) );
  NAND2X0 U302 ( .IN1(n206), .IN2(reg_a[21]), .QN(n482) );
  NAND2X1 U303 ( .IN1(n537), .IN2(n540), .QN(n360) );
  NOR2X4 U304 ( .IN1(n152), .IN2(n111), .QN(n178) );
  INVX0 U305 ( .IN(n354), .QN(n382) );
  OR2X1 U306 ( .IN1(reg_a[23]), .IN2(n343), .Q(n345) );
  INVX0 U307 ( .IN(n412), .QN(n414) );
  NOR2X0 U308 ( .IN1(n506), .IN2(n107), .QN(n394) );
  NAND2X0 U309 ( .IN1(n191), .IN2(n100), .QN(n413) );
  INVX0 U310 ( .IN(n229), .QN(n247) );
  NAND2X2 U311 ( .IN1(n428), .IN2(n109), .QN(n378) );
  NOR2X4 U312 ( .IN1(n379), .IN2(n378), .QN(n434) );
  OA21X1 U313 ( .IN1(n250), .IN2(n487), .IN3(n486), .Q(n488) );
  NAND2X0 U314 ( .IN1(n207), .IN2(reg_a[9]), .QN(n428) );
  OAI21X1 U315 ( .IN1(reg_a[22]), .IN2(n208), .IN3(n481), .QN(n487) );
  NOR2X4 U316 ( .IN1(n177), .IN2(n119), .QN(n152) );
  NOR2X4 U317 ( .IN1(n104), .IN2(n214), .QN(n148) );
  NOR2X4 U318 ( .IN1(n104), .IN2(n214), .QN(n149) );
  INVX0 U319 ( .IN(n104), .QN(n171) );
  INVX0 U320 ( .IN(n487), .QN(n175) );
  OR2X1 U321 ( .IN1(n116), .IN2(n140), .Q(n555) );
  NOR2X0 U322 ( .IN1(n253), .IN2(n478), .QN(n154) );
  AND2X1 U323 ( .IN1(n164), .IN2(reg_b[3]), .Q(n362) );
  NAND2X0 U324 ( .IN1(reg_b[31]), .IN2(n155), .QN(n409) );
  XOR3X1 U325 ( .IN1(n204), .IN2(reg_a[10]), .IN3(n156), .Q(n431) );
  OAI21X1 U326 ( .IN1(n429), .IN2(n181), .IN3(n428), .QN(n156) );
  XOR3X1 U327 ( .IN1(n157), .IN2(reg_a[16]), .IN3(n158), .Q(n459) );
  OAI21X1 U328 ( .IN1(n457), .IN2(n185), .IN3(n456), .QN(n158) );
  XOR3X1 U329 ( .IN1(reg_b[19]), .IN2(n159), .IN3(n160), .Q(n472) );
  OAI21X1 U330 ( .IN1(n470), .IN2(n183), .IN3(n469), .QN(n160) );
  XOR3X1 U331 ( .IN1(reg_b[20]), .IN2(n161), .IN3(n162), .Q(n477) );
  OAI21X1 U332 ( .IN1(n475), .IN2(n474), .IN3(n473), .QN(n162) );
  XOR3X1 U333 ( .IN1(n208), .IN2(reg_a[22]), .IN3(n163), .Q(n485) );
  OAI21X1 U334 ( .IN1(n483), .IN2(n154), .IN3(n482), .QN(n163) );
  OR2X1 U335 ( .IN1(n164), .IN2(reg_b[3]), .Q(n365) );
  NAND2X0 U336 ( .IN1(n223), .IN2(n222), .QN(n537) );
  OR2X1 U337 ( .IN1(reg_a[9]), .IN2(n207), .Q(n427) );
  OR2X1 U338 ( .IN1(reg_b[13]), .IN2(n165), .Q(n447) );
  OAI21X1 U339 ( .IN1(reg_a[10]), .IN2(n204), .IN3(n427), .QN(n433) );
  OR2X1 U340 ( .IN1(reg_a[8]), .IN2(n125), .Q(n376) );
  OR2X1 U341 ( .IN1(reg_b[16]), .IN2(n166), .Q(n460) );
  NAND2X0 U342 ( .IN1(reg_b[28]), .IN2(n190), .QN(n399) );
  NOR2X4 U343 ( .IN1(n434), .IN2(n121), .QN(n177) );
  NBUFFX2 U344 ( .IN(n581), .Q(n257) );
  NBUFFX2 U345 ( .IN(n581), .Q(n259) );
  NBUFFX2 U346 ( .IN(n581), .Q(n263) );
  NBUFFX2 U347 ( .IN(n581), .Q(n262) );
  NBUFFX2 U348 ( .IN(n581), .Q(n261) );
  NBUFFX2 U349 ( .IN(n581), .Q(n260) );
  NBUFFX2 U350 ( .IN(n581), .Q(n264) );
  INVX0 U351 ( .IN(n299), .QN(n289) );
  INVX0 U352 ( .IN(n298), .QN(n291) );
  INVX0 U353 ( .IN(n299), .QN(n290) );
  INVX0 U354 ( .IN(n298), .QN(n292) );
  INVX0 U355 ( .IN(n297), .QN(n294) );
  INVX0 U356 ( .IN(n296), .QN(n295) );
  INVX0 U357 ( .IN(n297), .QN(n293) );
  INVX0 U358 ( .IN(n275), .QN(n299) );
  INVX0 U359 ( .IN(n275), .QN(n298) );
  INVX0 U360 ( .IN(n6), .QN(n300) );
  INVX0 U361 ( .IN(n282), .QN(n301) );
  INVX0 U362 ( .IN(n276), .QN(n302) );
  INVX0 U363 ( .IN(n277), .QN(n304) );
  INVX0 U364 ( .IN(n277), .QN(n305) );
  INVX0 U365 ( .IN(n278), .QN(n306) );
  INVX0 U366 ( .IN(n278), .QN(n307) );
  INVX0 U367 ( .IN(n279), .QN(n308) );
  INVX0 U368 ( .IN(n279), .QN(n309) );
  INVX0 U369 ( .IN(n280), .QN(n310) );
  INVX0 U370 ( .IN(n280), .QN(n311) );
  INVX0 U371 ( .IN(n281), .QN(n312) );
  INVX0 U372 ( .IN(n276), .QN(n303) );
  INVX0 U373 ( .IN(n282), .QN(n315) );
  INVX0 U374 ( .IN(n281), .QN(n313) );
  INVX0 U375 ( .IN(n282), .QN(n314) );
  NOR2X0 U376 ( .IN1(n172), .IN2(n417), .QN(n169) );
  INVX0 U377 ( .IN(n555), .QN(n372) );
  OR2X1 U378 ( .IN1(n359), .IN2(n153), .Q(n416) );
  INVX0 U379 ( .IN(n274), .QN(n296) );
  INVX0 U380 ( .IN(n287), .QN(n275) );
  INVX0 U381 ( .IN(n286), .QN(n276) );
  INVX0 U382 ( .IN(n286), .QN(n277) );
  INVX0 U383 ( .IN(n274), .QN(n297) );
  INVX0 U384 ( .IN(n285), .QN(n278) );
  INVX0 U385 ( .IN(n285), .QN(n279) );
  INVX0 U386 ( .IN(n284), .QN(n280) );
  INVX0 U387 ( .IN(n284), .QN(n281) );
  INVX0 U388 ( .IN(n283), .QN(n282) );
  OR2X1 U389 ( .IN1(n529), .IN2(n522), .Q(n402) );
  NOR2X0 U390 ( .IN1(n124), .IN2(n416), .QN(n172) );
  NOR2X0 U391 ( .IN1(n172), .IN2(n551), .QN(n173) );
  INVX0 U392 ( .IN(n411), .QN(n245) );
  INVX0 U393 ( .IN(n411), .QN(n246) );
  OR2X1 U394 ( .IN1(n522), .IN2(n531), .Q(n525) );
  OR2X1 U395 ( .IN1(n529), .IN2(n561), .Q(n533) );
  INVX0 U396 ( .IN(n554), .QN(n556) );
  INVX0 U397 ( .IN(n469), .QN(n385) );
  INVX0 U398 ( .IN(n376), .QN(n368) );
  NOR2X0 U399 ( .IN1(n571), .IN2(n570), .QN(n575) );
  NOR2X0 U400 ( .IN1(n126), .IN2(n566), .QN(n571) );
  INVX0 U401 ( .IN(n456), .QN(n383) );
  INVX0 U402 ( .IN(n442), .QN(n381) );
  NOR2X0 U403 ( .IN1(n521), .IN2(n402), .QN(n404) );
  NOR2X0 U404 ( .IN1(n510), .IN2(n509), .QN(n515) );
  NOR2X0 U405 ( .IN1(n126), .IN2(n501), .QN(n510) );
  INVX0 U406 ( .IN(n482), .QN(n388) );
  INVX0 U407 ( .IN(n6), .QN(n287) );
  INVX0 U408 ( .IN(n6), .QN(n286) );
  INVX0 U409 ( .IN(n6), .QN(n285) );
  INVX0 U410 ( .IN(n6), .QN(n284) );
  INVX0 U411 ( .IN(n6), .QN(n283) );
  INVX0 U412 ( .IN(n288), .QN(n274) );
  INVX0 U413 ( .IN(n6), .QN(n288) );
  OR2X1 U414 ( .IN1(n584), .IN2(n210), .Q(n412) );
  OR3X1 U415 ( .IN1(n210), .IN2(n586), .IN3(n241), .Q(gcd_ns[0]) );
  AND2X1 U416 ( .IN1(n584), .IN2(n280), .Q(n586) );
  OA21X1 U417 ( .IN1(n169), .IN2(n424), .IN3(n109), .Q(n181) );
  INVX0 U418 ( .IN(n413), .QN(n584) );
  INVX0 U419 ( .IN(n502), .QN(n503) );
  INVX0 U420 ( .IN(n528), .QN(n561) );
  INVX0 U421 ( .IN(n521), .QN(n531) );
  INVX0 U422 ( .IN(n530), .QN(n522) );
  INVX0 U423 ( .IN(n560), .QN(n529) );
  NOR2X0 U424 ( .IN1(n492), .IN2(n491), .QN(n182) );
  NOR2X0 U425 ( .IN1(n150), .IN2(n465), .QN(n183) );
  NOR2X0 U426 ( .IN1(n177), .IN2(n438), .QN(n184) );
  NOR2X0 U427 ( .IN1(n147), .IN2(n452), .QN(n185) );
  INVX0 U428 ( .IN(n348), .QN(n387) );
  INVX0 U429 ( .IN(n539), .QN(n541) );
  INVX0 U430 ( .IN(n427), .QN(n429) );
  INVX0 U431 ( .IN(n455), .QN(n457) );
  INVX0 U432 ( .IN(n468), .QN(n470) );
  INVX0 U433 ( .IN(n481), .QN(n483) );
  INVX0 U434 ( .IN(n495), .QN(n497) );
  INVX0 U435 ( .IN(n441), .QN(n443) );
  NBUFFX2 U436 ( .IN(n334), .Q(n329) );
  NBUFFX2 U437 ( .IN(n333), .Q(n331) );
  NBUFFX2 U438 ( .IN(n335), .Q(n328) );
  NBUFFX2 U439 ( .IN(n340), .Q(n317) );
  NBUFFX2 U440 ( .IN(n340), .Q(n318) );
  NBUFFX2 U441 ( .IN(n339), .Q(n319) );
  NBUFFX2 U442 ( .IN(n339), .Q(n320) );
  NBUFFX2 U443 ( .IN(n338), .Q(n321) );
  NBUFFX2 U444 ( .IN(n338), .Q(n322) );
  NBUFFX2 U445 ( .IN(n337), .Q(n323) );
  NBUFFX2 U446 ( .IN(n337), .Q(n324) );
  NBUFFX2 U447 ( .IN(n336), .Q(n325) );
  NBUFFX2 U448 ( .IN(n336), .Q(n326) );
  NBUFFX2 U449 ( .IN(n335), .Q(n327) );
  NBUFFX2 U450 ( .IN(n334), .Q(n330) );
  NBUFFX2 U451 ( .IN(n333), .Q(n332) );
  INVX0 U452 ( .IN(n418), .QN(n377) );
  AO222X1 U453 ( .IN1(n247), .IN2(reg_a[31]), .IN3(b_in[31]), .IN4(n102), 
        .IN5(reg_b[31]), .IN6(n256), .Q(N123) );
  AO222X1 U454 ( .IN1(n232), .IN2(reg_a[20]), .IN3(b_in[20]), .IN4(n102), 
        .IN5(reg_b[20]), .IN6(n256), .Q(N112) );
  AO222X1 U455 ( .IN1(n230), .IN2(reg_a[22]), .IN3(b_in[22]), .IN4(n170), 
        .IN5(reg_b[22]), .IN6(n256), .Q(N114) );
  AO222X1 U456 ( .IN1(n246), .IN2(reg_a[23]), .IN3(b_in[23]), .IN4(n102), 
        .IN5(reg_b[23]), .IN6(n255), .Q(N115) );
  AO222X1 U457 ( .IN1(n248), .IN2(reg_a[10]), .IN3(b_in[10]), .IN4(n170), 
        .IN5(reg_b[10]), .IN6(n255), .Q(N102) );
  AO222X1 U458 ( .IN1(n239), .IN2(reg_a[11]), .IN3(b_in[11]), .IN4(n170), 
        .IN5(reg_b[11]), .IN6(n255), .Q(N103) );
  AO222X1 U459 ( .IN1(n235), .IN2(reg_a[14]), .IN3(b_in[14]), .IN4(n102), 
        .IN5(reg_b[14]), .IN6(n255), .Q(N106) );
  AO222X1 U460 ( .IN1(n247), .IN2(reg_a[15]), .IN3(b_in[15]), .IN4(n170), 
        .IN5(reg_b[15]), .IN6(n255), .Q(N107) );
  AO222X1 U461 ( .IN1(n245), .IN2(reg_a[16]), .IN3(b_in[16]), .IN4(n170), 
        .IN5(reg_b[16]), .IN6(n255), .Q(N108) );
  AO222X1 U462 ( .IN1(n248), .IN2(reg_a[17]), .IN3(b_in[17]), .IN4(n102), 
        .IN5(reg_b[17]), .IN6(n255), .Q(N109) );
  AO222X1 U463 ( .IN1(n233), .IN2(reg_a[25]), .IN3(b_in[25]), .IN4(n170), 
        .IN5(reg_b[25]), .IN6(n256), .Q(N117) );
  AO222X1 U464 ( .IN1(n238), .IN2(reg_a[27]), .IN3(b_in[27]), .IN4(n170), 
        .IN5(reg_b[27]), .IN6(n255), .Q(N119) );
  AO222X1 U465 ( .IN1(n237), .IN2(reg_a[29]), .IN3(b_in[29]), .IN4(n102), 
        .IN5(reg_b[29]), .IN6(n256), .Q(N121) );
  AO222X1 U466 ( .IN1(n232), .IN2(reg_a[3]), .IN3(b_in[3]), .IN4(n102), .IN5(
        reg_b[3]), .IN6(n255), .Q(N95) );
  NAND2X0 U467 ( .IN1(n187), .IN2(reg_b[2]), .QN(n539) );
  AND3X1 U468 ( .IN1(reg_a[31]), .IN2(n563), .IN3(n562), .Q(n565) );
  OAI21X1 U469 ( .IN1(n561), .IN2(n174), .IN3(n560), .QN(n562) );
  MUX21X1 U470 ( .IN1(n525), .IN2(n524), .S(n110), .Q(n527) );
  XOR2X1 U471 ( .IN1(n201), .IN2(reg_a[29]), .Q(n524) );
  XOR3X1 U472 ( .IN1(n211), .IN2(n106), .IN3(n548), .Q(n550) );
  XOR3X1 U473 ( .IN1(reg_b[3]), .IN2(reg_a[3]), .IN3(n542), .Q(n544) );
  OA21X1 U474 ( .IN1(n541), .IN2(n180), .IN3(n540), .Q(n542) );
  XOR3X1 U475 ( .IN1(n216), .IN2(n116), .IN3(n173), .Q(n553) );
  XOR3X1 U476 ( .IN1(reg_b[25]), .IN2(reg_a[25]), .IN3(n498), .Q(n500) );
  OA21X1 U477 ( .IN1(n497), .IN2(n182), .IN3(n496), .Q(n498) );
  XOR3X1 U478 ( .IN1(reg_b[14]), .IN2(reg_a[14]), .IN3(n449), .Q(n451) );
  XOR3X1 U479 ( .IN1(reg_b[23]), .IN2(reg_a[23]), .IN3(n488), .Q(n490) );
  XOR3X1 U480 ( .IN1(reg_b[8]), .IN2(reg_a[8]), .IN3(n420), .Q(n423) );
  AND2X1 U481 ( .IN1(reg_b[1]), .IN2(n128), .Q(n572) );
  AND2X1 U482 ( .IN1(reg_b[26]), .IN2(n148), .Q(n512) );
  XOR3X1 U483 ( .IN1(reg_b[28]), .IN2(reg_a[28]), .IN3(n122), .Q(n520) );
  MUX21X1 U484 ( .IN1(n533), .IN2(n532), .S(n174), .Q(n535) );
  XOR2X1 U485 ( .IN1(n202), .IN2(reg_a[30]), .Q(n532) );
  XOR3X1 U486 ( .IN1(reg_a[12]), .IN2(reg_b[12]), .IN3(n184), .Q(n440) );
  XOR3X1 U487 ( .IN1(reg_a[15]), .IN2(reg_b[15]), .IN3(n185), .Q(n454) );
  XOR3X1 U488 ( .IN1(reg_a[9]), .IN2(reg_b[9]), .IN3(n181), .Q(n426) );
  XOR3X1 U489 ( .IN1(reg_a[18]), .IN2(reg_b[18]), .IN3(n183), .Q(n467) );
  XOR3X1 U490 ( .IN1(reg_a[21]), .IN2(reg_b[21]), .IN3(n154), .Q(n480) );
  XOR3X1 U491 ( .IN1(reg_a[24]), .IN2(reg_b[24]), .IN3(n182), .Q(n494) );
  OA21X1 U492 ( .IN1(n443), .IN2(n184), .IN3(n442), .Q(n444) );
  OA21X1 U493 ( .IN1(n556), .IN2(n173), .IN3(n555), .Q(n557) );
  XOR3X1 U494 ( .IN1(reg_b[11]), .IN2(reg_a[11]), .IN3(n435), .Q(n437) );
  XOR3X1 U495 ( .IN1(reg_b[17]), .IN2(reg_a[17]), .IN3(n462), .Q(n464) );
  OAI21X1 U496 ( .IN1(reg_b[0]), .IN2(n578), .IN3(n577), .QN(n582) );
  INVX0 U497 ( .IN(reg_a[0]), .QN(n578) );
  XOR3X1 U498 ( .IN1(reg_b[26]), .IN2(reg_a[26]), .IN3(n507), .Q(n508) );
  OAI21X1 U499 ( .IN1(reg_a[25]), .IN2(n205), .IN3(n495), .QN(n502) );
  AO22X1 U500 ( .IN1(n344), .IN2(n345), .IN3(reg_a[23]), .IN4(n343), .Q(n491)
         );
  AO22X1 U501 ( .IN1(n353), .IN2(n354), .IN3(reg_a[14]), .IN4(n352), .Q(n452)
         );
  INVX0 U502 ( .IN(n447), .QN(n353) );
  AO22X1 U503 ( .IN1(n357), .IN2(n358), .IN3(reg_a[11]), .IN4(n356), .Q(n438)
         );
  INVX0 U504 ( .IN(n432), .QN(n357) );
  OR4X1 U505 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n63) );
  OR4X1 U506 ( .IN1(n116), .IN2(reg_b[7]), .IN3(reg_b[8]), .IN4(reg_b[9]), .Q(
        n59) );
  OR4X1 U507 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n62) );
  OR4X1 U508 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(
        reg_b[16]), .Q(n65) );
  OR2X1 U509 ( .IN1(reg_a[30]), .IN2(n202), .Q(n528) );
  OR2X1 U510 ( .IN1(reg_a[29]), .IN2(n201), .Q(n521) );
  AO22X1 U511 ( .IN1(reg_a[8]), .IN2(n300), .IN3(result[8]), .IN4(n276), .Q(
        n68) );
  AO22X1 U512 ( .IN1(reg_a[9]), .IN2(n301), .IN3(result[9]), .IN4(n295), .Q(
        n69) );
  AO22X1 U513 ( .IN1(reg_a[10]), .IN2(n301), .IN3(result[10]), .IN4(n295), .Q(
        n70) );
  AO22X1 U514 ( .IN1(reg_a[11]), .IN2(n302), .IN3(result[11]), .IN4(n295), .Q(
        n71) );
  AO22X1 U515 ( .IN1(reg_a[12]), .IN2(n302), .IN3(result[12]), .IN4(n295), .Q(
        n72) );
  AO22X1 U516 ( .IN1(reg_a[14]), .IN2(n303), .IN3(result[14]), .IN4(n294), .Q(
        n74) );
  AO22X1 U517 ( .IN1(reg_a[15]), .IN2(n304), .IN3(result[15]), .IN4(n294), .Q(
        n75) );
  AO22X1 U518 ( .IN1(reg_a[16]), .IN2(n304), .IN3(result[16]), .IN4(n294), .Q(
        n76) );
  AO22X1 U519 ( .IN1(reg_a[17]), .IN2(n305), .IN3(result[17]), .IN4(n293), .Q(
        n77) );
  AO22X1 U520 ( .IN1(reg_a[18]), .IN2(n305), .IN3(result[18]), .IN4(n293), .Q(
        n78) );
  AO22X1 U521 ( .IN1(reg_a[19]), .IN2(n306), .IN3(result[19]), .IN4(n293), .Q(
        n79) );
  AO22X1 U522 ( .IN1(reg_a[20]), .IN2(n306), .IN3(result[20]), .IN4(n293), .Q(
        n80) );
  AO22X1 U523 ( .IN1(reg_a[21]), .IN2(n307), .IN3(result[21]), .IN4(n292), .Q(
        n81) );
  AO22X1 U524 ( .IN1(reg_a[22]), .IN2(n307), .IN3(result[22]), .IN4(n292), .Q(
        n82) );
  AO22X1 U525 ( .IN1(reg_a[23]), .IN2(n308), .IN3(result[23]), .IN4(n292), .Q(
        n83) );
  AO22X1 U526 ( .IN1(reg_a[24]), .IN2(n308), .IN3(result[24]), .IN4(n291), .Q(
        n84) );
  AO22X1 U527 ( .IN1(reg_a[25]), .IN2(n309), .IN3(result[25]), .IN4(n291), .Q(
        n85) );
  AO22X1 U528 ( .IN1(reg_a[26]), .IN2(n309), .IN3(result[26]), .IN4(n291), .Q(
        n86) );
  AO22X1 U529 ( .IN1(reg_a[27]), .IN2(n310), .IN3(result[27]), .IN4(n291), .Q(
        n87) );
  AO22X1 U530 ( .IN1(reg_a[28]), .IN2(n310), .IN3(result[28]), .IN4(n290), .Q(
        n88) );
  AO22X1 U531 ( .IN1(reg_a[29]), .IN2(n311), .IN3(result[29]), .IN4(n290), .Q(
        n89) );
  AO22X1 U532 ( .IN1(reg_a[30]), .IN2(n311), .IN3(result[30]), .IN4(n290), .Q(
        n90) );
  AO22X1 U533 ( .IN1(reg_a[2]), .IN2(n312), .IN3(result[2]), .IN4(n290), .Q(
        n91) );
  AO22X1 U534 ( .IN1(reg_a[3]), .IN2(n312), .IN3(result[3]), .IN4(n289), .Q(
        n92) );
  AO22X1 U535 ( .IN1(reg_a[31]), .IN2(n315), .IN3(result[31]), .IN4(n278), .Q(
        n97) );
  AO22X1 U536 ( .IN1(reg_a[0]), .IN2(n301), .IN3(result[0]), .IN4(n292), .Q(
        n99) );
  NAND2X0 U537 ( .IN1(n196), .IN2(reg_a[24]), .QN(n496) );
  NAND2X0 U538 ( .IN1(n201), .IN2(reg_a[29]), .QN(n530) );
  NAND2X0 U539 ( .IN1(n202), .IN2(reg_a[30]), .QN(n560) );
  NAND2X0 U540 ( .IN1(reg_a[26]), .IN2(n342), .QN(n392) );
  NAND2X0 U541 ( .IN1(reg_a[31]), .IN2(n563), .QN(n407) );
  NAND2X0 U542 ( .IN1(n205), .IN2(reg_a[25]), .QN(n506) );
  NAND2X0 U543 ( .IN1(reg_b[27]), .IN2(n398), .QN(n396) );
  OAI21X1 U544 ( .IN1(reg_a[16]), .IN2(n157), .IN3(n455), .QN(n461) );
  NAND2X0 U545 ( .IN1(n208), .IN2(reg_a[22]), .QN(n486) );
  AND2X1 U546 ( .IN1(n209), .IN2(n67), .Q(done) );
  AND3X1 U547 ( .IN1(start), .IN2(n67), .IN3(n100), .Q(n210) );
  AO22X1 U548 ( .IN1(n350), .IN2(n351), .IN3(reg_a[17]), .IN4(n349), .Q(n465)
         );
  NBUFFX2 U549 ( .IN(n341), .Q(n316) );
  NBUFFX2 U550 ( .IN(reset_n), .Q(n341) );
  INVX0 U551 ( .IN(a_in[1]), .QN(n566) );
  INVX0 U552 ( .IN(a_in[26]), .QN(n501) );
  NBUFFX2 U553 ( .IN(reset_n), .Q(n340) );
  NBUFFX2 U554 ( .IN(reset_n), .Q(n339) );
  NBUFFX2 U555 ( .IN(reset_n), .Q(n338) );
  NBUFFX2 U556 ( .IN(reset_n), .Q(n337) );
  NBUFFX2 U557 ( .IN(reset_n), .Q(n336) );
  NBUFFX2 U558 ( .IN(reset_n), .Q(n335) );
  NBUFFX2 U559 ( .IN(reset_n), .Q(n334) );
  NBUFFX2 U560 ( .IN(reset_n), .Q(n333) );
  XOR3X1 U561 ( .IN1(reg_b[13]), .IN2(reg_a[13]), .IN3(n444), .Q(n446) );
  OAI21X1 U562 ( .IN1(reg_a[13]), .IN2(n355), .IN3(n441), .QN(n448) );
  AO22X1 U563 ( .IN1(reg_a[13]), .IN2(n303), .IN3(result[13]), .IN4(n294), .Q(
        n73) );
  AO222X1 U564 ( .IN1(n247), .IN2(reg_a[7]), .IN3(b_in[7]), .IN4(n170), .IN5(
        reg_b[7]), .IN6(n256), .Q(N99) );
  XOR3X1 U565 ( .IN1(reg_b[7]), .IN2(reg_a[7]), .IN3(n557), .Q(n559) );
  AO22X1 U566 ( .IN1(reg_a[7]), .IN2(n314), .IN3(result[7]), .IN4(n281), .Q(
        n96) );
  INVX8 U567 ( .IN(n141), .QN(n212) );
  INVX8 U568 ( .IN(n141), .QN(n213) );
  INVX8 U569 ( .IN(n141), .QN(n579) );
  AO22X1 U570 ( .IN1(n222), .IN2(n315), .IN3(result[1]), .IN4(n279), .Q(n98)
         );
  OA21X1 U571 ( .IN1(n169), .IN2(n419), .IN3(n418), .Q(n420) );
  OA21X1 U572 ( .IN1(n124), .IN2(n153), .IN3(n547), .Q(n548) );
  NOR2X0 U573 ( .IN1(n569), .IN2(n568), .QN(n570) );
  NOR2X0 U574 ( .IN1(n508), .IN2(n568), .QN(n509) );
  AO222X1 U575 ( .IN1(n230), .IN2(reg_a[2]), .IN3(b_in[2]), .IN4(n102), .IN5(
        reg_b[2]), .IN6(n256), .Q(N94) );
  OR4X1 U576 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n61) );
  AO221X1 U577 ( .IN1(n583), .IN2(n485), .IN3(a_in[22]), .IN4(n260), .IN5(n484), .Q(N81) );
  NBUFFX2 U578 ( .IN(n265), .Q(n244) );
  AO222X1 U579 ( .IN1(n236), .IN2(reg_a[30]), .IN3(b_in[30]), .IN4(n170), 
        .IN5(reg_b[30]), .IN6(n255), .Q(N122) );
  NBUFFX2 U580 ( .IN(n271), .Q(n236) );
  AO222X1 U581 ( .IN1(n234), .IN2(reg_a[24]), .IN3(b_in[24]), .IN4(n102), 
        .IN5(reg_b[24]), .IN6(n255), .Q(N116) );
  NBUFFX2 U582 ( .IN(n272), .Q(n234) );
  AO222X1 U583 ( .IN1(n240), .IN2(reg_a[19]), .IN3(b_in[19]), .IN4(n170), 
        .IN5(reg_b[19]), .IN6(n255), .Q(N111) );
  NBUFFX2 U584 ( .IN(n268), .Q(n240) );
  AO222X1 U585 ( .IN1(n243), .IN2(reg_a[12]), .IN3(b_in[12]), .IN4(n170), 
        .IN5(reg_b[12]), .IN6(n255), .Q(N104) );
  NBUFFX2 U586 ( .IN(n266), .Q(n243) );
  OR4X1 U587 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(
        reg_b[1]), .Q(n64) );
  NAND2X0 U588 ( .IN1(n504), .IN2(n503), .QN(n505) );
  AO22X1 U589 ( .IN1(n371), .IN2(n370), .IN3(n211), .IN4(n220), .Q(n551) );
  AO22X1 U590 ( .IN1(n211), .IN2(n313), .IN3(result[5]), .IN4(n289), .Q(n94)
         );
  AO222X1 U591 ( .IN1(n242), .IN2(n216), .IN3(b_in[6]), .IN4(n170), .IN5(n116), 
        .IN6(n256), .Q(N98) );
  AO22X1 U592 ( .IN1(n216), .IN2(n314), .IN3(result[6]), .IN4(n289), .Q(n95)
         );
  OR4X1 U593 ( .IN1(reg_b[31]), .IN2(reg_b[3]), .IN3(n105), .IN4(n106), .Q(n60) );
  AO222X1 U594 ( .IN1(n231), .IN2(n221), .IN3(b_in[4]), .IN4(n170), .IN5(n105), 
        .IN6(n255), .Q(N96) );
  XOR3X1 U595 ( .IN1(n221), .IN2(n105), .IN3(n124), .Q(n546) );
  AO22X1 U596 ( .IN1(n221), .IN2(n313), .IN3(result[4]), .IN4(n289), .Q(n93)
         );
  INVX2 U597 ( .IN(n224), .QN(n225) );
  AO221X1 U598 ( .IN1(n130), .IN2(n464), .IN3(a_in[17]), .IN4(n262), .IN5(n463), .Q(N76) );
  AO222X1 U599 ( .IN1(n245), .IN2(reg_a[9]), .IN3(b_in[9]), .IN4(n170), .IN5(
        reg_b[9]), .IN6(n255), .Q(N101) );
  AO222X1 U600 ( .IN1(n231), .IN2(reg_a[21]), .IN3(b_in[21]), .IN4(n102), 
        .IN5(reg_b[21]), .IN6(n256), .Q(N113) );
  AO222X1 U601 ( .IN1(n247), .IN2(reg_a[18]), .IN3(b_in[18]), .IN4(n102), 
        .IN5(reg_b[18]), .IN6(n256), .Q(N110) );
  AO222X1 U602 ( .IN1(n245), .IN2(reg_a[28]), .IN3(b_in[28]), .IN4(n170), 
        .IN5(reg_b[28]), .IN6(n256), .Q(N120) );
  AO222X1 U603 ( .IN1(n267), .IN2(n211), .IN3(b_in[5]), .IN4(n102), .IN5(n106), 
        .IN6(n256), .Q(N97) );
  AO222X1 U604 ( .IN1(n246), .IN2(n222), .IN3(b_in[1]), .IN4(n102), .IN5(
        reg_b[1]), .IN6(n255), .Q(N93) );
  AO222X1 U605 ( .IN1(n248), .IN2(reg_a[26]), .IN3(b_in[26]), .IN4(n170), 
        .IN5(reg_b[26]), .IN6(n256), .Q(N118) );
  AO222X1 U606 ( .IN1(n246), .IN2(reg_a[13]), .IN3(b_in[13]), .IN4(n102), 
        .IN5(reg_b[13]), .IN6(n256), .Q(N105) );
  AO222X1 U607 ( .IN1(n244), .IN2(reg_a[8]), .IN3(b_in[8]), .IN4(n102), .IN5(
        reg_b[8]), .IN6(n256), .Q(N100) );
  NOR2X0 U608 ( .IN1(n146), .IN2(n219), .QN(n573) );
  NOR2X0 U609 ( .IN1(n511), .IN2(n219), .QN(n513) );
  AO221X1 U610 ( .IN1(n583), .IN2(n446), .IN3(a_in[13]), .IN4(n263), .IN5(n445), .Q(N72) );
  NBUFFX2 U611 ( .IN(n585), .Q(n230) );
  NBUFFX2 U612 ( .IN(n585), .Q(n231) );
  NBUFFX2 U613 ( .IN(n273), .Q(n232) );
  NBUFFX2 U614 ( .IN(n272), .Q(n233) );
  NBUFFX2 U615 ( .IN(n271), .Q(n235) );
  NBUFFX2 U616 ( .IN(n270), .Q(n237) );
  NBUFFX2 U617 ( .IN(n269), .Q(n238) );
  NBUFFX2 U618 ( .IN(n268), .Q(n239) );
  NBUFFX2 U619 ( .IN(n267), .Q(n241) );
  NBUFFX2 U620 ( .IN(n266), .Q(n242) );
  NBUFFX2 U621 ( .IN(n585), .Q(n272) );
  NBUFFX2 U622 ( .IN(n585), .Q(n271) );
  NBUFFX2 U623 ( .IN(n585), .Q(n270) );
  NBUFFX2 U624 ( .IN(n585), .Q(n269) );
  NBUFFX2 U625 ( .IN(n585), .Q(n268) );
  NBUFFX2 U626 ( .IN(n585), .Q(n267) );
  NBUFFX2 U627 ( .IN(n585), .Q(n266) );
  NBUFFX2 U628 ( .IN(n585), .Q(n265) );
  AND3X1 U629 ( .IN1(n348), .IN2(n251), .IN3(n386), .Q(n249) );
  NOR3X0 U630 ( .IN1(n249), .IN2(n478), .IN3(n388), .QN(n250) );
  NOR3X0 U631 ( .IN1(n387), .IN2(n474), .IN3(n475), .QN(n253) );
  AO221X1 U632 ( .IN1(n130), .IN2(n459), .IN3(a_in[16]), .IN4(n262), .IN5(n458), .Q(N75) );
  AO221X1 U633 ( .IN1(n130), .IN2(n520), .IN3(a_in[28]), .IN4(n259), .IN5(n519), .Q(N87) );
  AO221X1 U634 ( .IN1(n130), .IN2(n544), .IN3(a_in[3]), .IN4(n258), .IN5(n543), 
        .Q(N62) );
  AO22X1 U635 ( .IN1(n149), .IN2(reg_b[12]), .IN3(n212), .IN4(reg_a[12]), .Q(
        n439) );
  AO221X1 U636 ( .IN1(n583), .IN2(n477), .IN3(a_in[20]), .IN4(n261), .IN5(n476), .Q(N79) );
  AO22X1 U637 ( .IN1(n128), .IN2(reg_b[20]), .IN3(n579), .IN4(reg_a[20]), .Q(
        n476) );
  AO221X1 U638 ( .IN1(n130), .IN2(n451), .IN3(a_in[14]), .IN4(n262), .IN5(n450), .Q(N73) );
  AO22X1 U639 ( .IN1(n149), .IN2(reg_b[14]), .IN3(n213), .IN4(reg_a[14]), .Q(
        n450) );
  AO221X1 U640 ( .IN1(n583), .IN2(n437), .IN3(a_in[11]), .IN4(n263), .IN5(n436), .Q(N70) );
  AO22X1 U641 ( .IN1(n149), .IN2(reg_b[11]), .IN3(n579), .IN4(reg_a[11]), .Q(
        n436) );
  AO221X1 U642 ( .IN1(n130), .IN2(n472), .IN3(a_in[19]), .IN4(n261), .IN5(n471), .Q(N78) );
  AO22X1 U643 ( .IN1(n148), .IN2(reg_b[19]), .IN3(n579), .IN4(reg_a[19]), .Q(
        n471) );
  AO221X1 U644 ( .IN1(n130), .IN2(n480), .IN3(a_in[21]), .IN4(n261), .IN5(n479), .Q(N80) );
  AO22X1 U645 ( .IN1(n149), .IN2(reg_b[21]), .IN3(n213), .IN4(reg_a[21]), .Q(
        n479) );
  AO221X1 U646 ( .IN1(n130), .IN2(n467), .IN3(a_in[18]), .IN4(n261), .IN5(n466), .Q(N77) );
  AO22X1 U647 ( .IN1(n128), .IN2(reg_b[18]), .IN3(n579), .IN4(reg_a[18]), .Q(
        n466) );
  AO221X1 U648 ( .IN1(n130), .IN2(n454), .IN3(a_in[15]), .IN4(n262), .IN5(n453), .Q(N74) );
  AO22X1 U649 ( .IN1(n149), .IN2(reg_b[15]), .IN3(n212), .IN4(reg_a[15]), .Q(
        n453) );
  AO22X1 U650 ( .IN1(n148), .IN2(reg_b[0]), .IN3(n213), .IN4(reg_a[0]), .Q(
        n580) );
  AO22X1 U651 ( .IN1(n148), .IN2(reg_b[13]), .IN3(n213), .IN4(reg_a[13]), .Q(
        n445) );
  AO221X1 U652 ( .IN1(n583), .IN2(n431), .IN3(a_in[10]), .IN4(n263), .IN5(n430), .Q(N69) );
  AO22X1 U653 ( .IN1(n149), .IN2(reg_b[10]), .IN3(n212), .IN4(reg_a[10]), .Q(
        n430) );
  AO22X1 U654 ( .IN1(n149), .IN2(n105), .IN3(n579), .IN4(n221), .Q(n545) );
  OA21X1 U655 ( .IN1(n151), .IN2(n461), .IN3(n460), .Q(n462) );
  AO221X1 U656 ( .IN1(n130), .IN2(n546), .IN3(a_in[4]), .IN4(n258), .IN5(n545), 
        .Q(N63) );
  AO22X1 U657 ( .IN1(n149), .IN2(reg_b[31]), .IN3(n579), .IN4(reg_a[31]), .Q(
        n564) );
  AO221X1 U658 ( .IN1(n130), .IN2(n423), .IN3(a_in[8]), .IN4(n264), .IN5(n422), 
        .Q(N67) );
  AO22X1 U659 ( .IN1(n148), .IN2(reg_b[8]), .IN3(n212), .IN4(reg_a[8]), .Q(
        n422) );
  AO221X1 U660 ( .IN1(n583), .IN2(n518), .IN3(a_in[27]), .IN4(n259), .IN5(n517), .Q(N86) );
  AO22X1 U661 ( .IN1(n149), .IN2(reg_b[27]), .IN3(n212), .IN4(reg_a[27]), .Q(
        n517) );
  AO221X1 U662 ( .IN1(n583), .IN2(n527), .IN3(a_in[29]), .IN4(n259), .IN5(n526), .Q(N88) );
  AO22X1 U663 ( .IN1(n148), .IN2(reg_b[29]), .IN3(n213), .IN4(reg_a[29]), .Q(
        n526) );
  AO221X1 U664 ( .IN1(n130), .IN2(n559), .IN3(a_in[7]), .IN4(n257), .IN5(n558), 
        .Q(N66) );
  AO22X1 U665 ( .IN1(n148), .IN2(reg_b[7]), .IN3(n579), .IN4(reg_a[7]), .Q(
        n558) );
  AO221X1 U666 ( .IN1(n583), .IN2(n500), .IN3(a_in[25]), .IN4(n260), .IN5(n499), .Q(N84) );
  AO22X1 U667 ( .IN1(n148), .IN2(reg_b[25]), .IN3(n212), .IN4(reg_a[25]), .Q(
        n499) );
  AO22X1 U668 ( .IN1(n128), .IN2(reg_b[16]), .IN3(n579), .IN4(reg_a[16]), .Q(
        n458) );
  AO22X1 U669 ( .IN1(n149), .IN2(reg_b[17]), .IN3(n212), .IN4(reg_a[17]), .Q(
        n463) );
  AO22X1 U670 ( .IN1(n128), .IN2(n106), .IN3(n213), .IN4(n211), .Q(n549) );
  OA21X1 U671 ( .IN1(n152), .IN2(n448), .IN3(n447), .Q(n449) );
  AO221X1 U672 ( .IN1(n583), .IN2(n490), .IN3(a_in[23]), .IN4(n260), .IN5(n489), .Q(N82) );
  AO22X1 U673 ( .IN1(n128), .IN2(reg_b[23]), .IN3(n213), .IN4(reg_a[23]), .Q(
        n489) );
  AO221X1 U674 ( .IN1(n583), .IN2(n550), .IN3(a_in[5]), .IN4(n258), .IN5(n549), 
        .Q(N64) );
  AO222X1 U675 ( .IN1(reg_a[0]), .IN2(n245), .IN3(b_in[0]), .IN4(n102), .IN5(
        reg_b[0]), .IN6(n256), .Q(N92) );
  OR4X1 U676 ( .IN1(reg_b[0]), .IN2(reg_b[10]), .IN3(reg_b[11]), .IN4(
        reg_b[12]), .Q(n66) );
  AO221X1 U677 ( .IN1(n583), .IN2(n535), .IN3(a_in[30]), .IN4(n259), .IN5(n534), .Q(N89) );
  AO22X1 U678 ( .IN1(n148), .IN2(reg_b[30]), .IN3(n213), .IN4(reg_a[30]), .Q(
        n534) );
  AO221X1 U679 ( .IN1(n130), .IN2(n553), .IN3(a_in[6]), .IN4(n257), .IN5(n552), 
        .Q(N65) );
  AO22X1 U680 ( .IN1(n128), .IN2(n116), .IN3(n212), .IN4(n216), .Q(n552) );
  AO221X1 U681 ( .IN1(n130), .IN2(n494), .IN3(a_in[24]), .IN4(n260), .IN5(n493), .Q(N83) );
  AO22X1 U682 ( .IN1(n128), .IN2(reg_b[24]), .IN3(n213), .IN4(reg_a[24]), .Q(
        n493) );
  AO22X1 U683 ( .IN1(n128), .IN2(reg_b[22]), .IN3(n579), .IN4(reg_a[22]), .Q(
        n484) );
  AO221X1 U684 ( .IN1(n130), .IN2(n426), .IN3(a_in[9]), .IN4(n264), .IN5(n425), 
        .Q(N68) );
  AO22X1 U685 ( .IN1(n148), .IN2(reg_b[9]), .IN3(n213), .IN4(reg_a[9]), .Q(
        n425) );
  AO221X1 U686 ( .IN1(n583), .IN2(n440), .IN3(a_in[12]), .IN4(n263), .IN5(n439), .Q(N71) );
  OA21X1 U687 ( .IN1(n434), .IN2(n433), .IN3(n432), .Q(n435) );
  AO221X1 U688 ( .IN1(n583), .IN2(n582), .IN3(a_in[0]), .IN4(n257), .IN5(n580), 
        .Q(N59) );
  AO221X1 U689 ( .IN1(n565), .IN2(n583), .IN3(a_in[31]), .IN4(n257), .IN5(n564), .Q(N90) );
  AO22X1 U690 ( .IN1(n128), .IN2(reg_b[28]), .IN3(n212), .IN4(reg_a[28]), .Q(
        n519) );
  NBUFFX2 U691 ( .IN(n585), .Q(n273) );
  AO22X1 U692 ( .IN1(n128), .IN2(reg_b[3]), .IN3(n212), .IN4(reg_a[3]), .Q(
        n543) );
  INVX4 U693 ( .IN(n516), .QN(n395) );
  OR2X2 U694 ( .IN1(n225), .IN2(n252), .Q(n577) );
  NAND2X4 U695 ( .IN1(n392), .IN2(n391), .QN(n393) );
  NOR2X4 U696 ( .IN1(n393), .IN2(n394), .QN(n516) );
  NAND2X4 U697 ( .IN1(n395), .IN2(n396), .QN(n397) );
  NAND2X4 U698 ( .IN1(n145), .IN2(n399), .QN(n400) );
  NAND2X4 U699 ( .IN1(n400), .IN2(n401), .QN(n523) );
  NOR2X4 U700 ( .IN1(n523), .IN2(n402), .QN(n403) );
  NOR2X4 U701 ( .IN1(n403), .IN2(n404), .QN(n405) );
  NAND2X4 U702 ( .IN1(n405), .IN2(n528), .QN(n406) );
  NAND2X4 U703 ( .IN1(n406), .IN2(n407), .QN(n408) );
  NAND2X4 U704 ( .IN1(n408), .IN2(n409), .QN(n410) );
endmodule

