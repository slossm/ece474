
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, n6, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ns;

  DFFARX1 \reg_b_reg[0]  ( .D(N92), .CLK(clk), .RSTB(n359), .Q(reg_b[0]), .QN(
        n273) );
  DFFARX1 \reg_b_reg[6]  ( .D(N98), .CLK(clk), .RSTB(n357), .Q(n113), .QN(n236) );
  DFFARX1 \reg_a_reg[4]  ( .D(N63), .CLK(clk), .RSTB(n356), .QN(n238) );
  DFFARX1 \reg_b_reg[1]  ( .D(N93), .CLK(clk), .RSTB(n359), .Q(reg_b[1]), .QN(
        n243) );
  DFFARX1 \reg_b_reg[4]  ( .D(N96), .CLK(clk), .RSTB(n356), .Q(n109), .QN(n152) );
  DFFARX1 \reg_a_reg[5]  ( .D(N64), .CLK(clk), .RSTB(n357), .QN(n156) );
  DFFARX1 \gcd_ps_reg[0]  ( .D(gcd_ns[0]), .CLK(clk), .RSTB(n360), .Q(n212), 
        .QN(n67) );
  DFFARX1 \reg_a_reg[20]  ( .D(N79), .CLK(clk), .RSTB(n350), .Q(reg_a[20]), 
        .QN(n180) );
  DFFARX1 \gcd_ps_reg[1]  ( .D(gcd_ns[1]), .CLK(clk), .RSTB(n359), .Q(n230), 
        .QN(n100) );
  DFFARX1 \reg_a_reg[13]  ( .D(N72), .CLK(clk), .RSTB(n346), .Q(reg_a[13]), 
        .QN(n184) );
  DFFARX1 \reg_b_reg[29]  ( .D(N121), .CLK(clk), .RSTB(n354), .Q(reg_b[29]), 
        .QN(n222) );
  DFFARX1 \reg_b_reg[30]  ( .D(N122), .CLK(clk), .RSTB(n355), .Q(reg_b[30]), 
        .QN(n223) );
  DFFARX1 \reg_a_reg[3]  ( .D(N62), .CLK(clk), .RSTB(n356), .Q(reg_a[3]), .QN(
        n183) );
  DFFARX1 \reg_a_reg[19]  ( .D(N78), .CLK(clk), .RSTB(n349), .Q(reg_a[19]), 
        .QN(n178) );
  DFFARX1 \reg_a_reg[16]  ( .D(N75), .CLK(clk), .RSTB(n348), .Q(reg_a[16]), 
        .QN(n185) );
  DFFARX1 \reg_a_reg[21]  ( .D(N80), .CLK(clk), .RSTB(n350), .Q(reg_a[21]), 
        .QN(n221) );
  DFFARX1 \reg_a_reg[12]  ( .D(N71), .CLK(clk), .RSTB(n346), .Q(reg_a[12]), 
        .QN(n224) );
  DFFARX1 \reg_a_reg[18]  ( .D(N77), .CLK(clk), .RSTB(n349), .Q(reg_a[18]), 
        .QN(n219) );
  DFFARX1 \reg_a_reg[24]  ( .D(N83), .CLK(clk), .RSTB(n352), .Q(reg_a[24]), 
        .QN(n218) );
  DFFARX1 \reg_a_reg[15]  ( .D(N74), .CLK(clk), .RSTB(n347), .Q(reg_a[15]), 
        .QN(n220) );
  DFFARX1 \reg_b_reg[25]  ( .D(N117), .CLK(clk), .RSTB(n352), .Q(reg_b[25]), 
        .QN(n226) );
  DFFARX1 \reg_b_reg[21]  ( .D(N113), .CLK(clk), .RSTB(n350), .Q(reg_b[21]), 
        .QN(n227) );
  DFFARX1 \reg_b_reg[10]  ( .D(N102), .CLK(clk), .RSTB(n345), .Q(reg_b[10]), 
        .QN(n225) );
  DFFARX1 \reg_b_reg[18]  ( .D(N110), .CLK(clk), .RSTB(n349), .Q(reg_b[18]), 
        .QN(n214) );
  DFFARX1 \reg_b_reg[22]  ( .D(N114), .CLK(clk), .RSTB(n351), .Q(reg_b[22]), 
        .QN(n229) );
  DFFARX1 \reg_b_reg[24]  ( .D(N116), .CLK(clk), .RSTB(n352), .Q(reg_b[24]), 
        .QN(n217) );
  DFFARX1 \reg_b_reg[19]  ( .D(N111), .CLK(clk), .RSTB(n349), .Q(reg_b[19]), 
        .QN(n216) );
  DFFARX1 \reg_b_reg[15]  ( .D(N107), .CLK(clk), .RSTB(n347), .Q(reg_b[15]), 
        .QN(n213) );
  DFFARX1 \reg_b_reg[16]  ( .D(N108), .CLK(clk), .RSTB(n348), .Q(reg_b[16]), 
        .QN(n176) );
  DFFARX1 \reg_b_reg[9]  ( .D(N101), .CLK(clk), .RSTB(n344), .Q(reg_b[9]), 
        .QN(n228) );
  DFFARX1 \reg_b_reg[12]  ( .D(N104), .CLK(clk), .RSTB(n346), .Q(reg_b[12]), 
        .QN(n215) );
  DFFARX1 \reg_a_reg[28]  ( .D(N87), .CLK(clk), .RSTB(n354), .Q(reg_a[28]), 
        .QN(n211) );
  DFFARX1 \reg_a_reg[31]  ( .D(N90), .CLK(clk), .RSTB(n358), .Q(reg_a[31]), 
        .QN(n174) );
  DFFARX1 \reg_a_reg[0]  ( .D(N59), .CLK(clk), .RSTB(n360), .Q(reg_a[0]), .QN(
        n244) );
  DFFARX1 \reg_a_reg[8]  ( .D(N67), .CLK(clk), .RSTB(n344), .QN(n129) );
  DFFARX1 \reg_b_reg[2]  ( .D(N94), .CLK(clk), .RSTB(n355), .Q(reg_b[2]), .QN(
        n210) );
  DFFARX1 \reg_b_reg[8]  ( .D(N100), .CLK(clk), .RSTB(n344), .Q(n106), .QN(
        n130) );
  DFFARX1 \reg_b_reg[7]  ( .D(N99), .CLK(clk), .RSTB(n358), .Q(n112), .QN(n209) );
  DFFARX1 \reg_a_reg[2]  ( .D(N61), .CLK(clk), .RSTB(n355), .QN(n208) );
  DFFARX1 \result_reg[31]  ( .D(n97), .CLK(clk), .RSTB(n358), .Q(result[31])
         );
  DFFARX1 \result_reg[7]  ( .D(n96), .CLK(clk), .RSTB(n358), .Q(result[7]) );
  DFFARX1 \result_reg[1]  ( .D(n98), .CLK(clk), .RSTB(n359), .Q(result[1]) );
  DFFARX1 \result_reg[8]  ( .D(n68), .CLK(clk), .RSTB(n344), .Q(result[8]) );
  DFFARX1 \result_reg[20]  ( .D(n80), .CLK(clk), .RSTB(n350), .Q(result[20])
         );
  DFFARX1 \result_reg[19]  ( .D(n79), .CLK(clk), .RSTB(n349), .Q(result[19])
         );
  DFFARX1 \result_reg[18]  ( .D(n78), .CLK(clk), .RSTB(n349), .Q(result[18])
         );
  DFFARX1 \result_reg[17]  ( .D(n77), .CLK(clk), .RSTB(n348), .Q(result[17])
         );
  DFFARX1 \result_reg[16]  ( .D(n76), .CLK(clk), .RSTB(n348), .Q(result[16])
         );
  DFFARX1 \result_reg[15]  ( .D(n75), .CLK(clk), .RSTB(n347), .Q(result[15])
         );
  DFFARX1 \result_reg[14]  ( .D(n74), .CLK(clk), .RSTB(n347), .Q(result[14])
         );
  DFFARX1 \result_reg[13]  ( .D(n73), .CLK(clk), .RSTB(n346), .Q(result[13])
         );
  DFFARX1 \result_reg[12]  ( .D(n72), .CLK(clk), .RSTB(n346), .Q(result[12])
         );
  DFFARX1 \result_reg[11]  ( .D(n71), .CLK(clk), .RSTB(n345), .Q(result[11])
         );
  DFFARX1 \result_reg[10]  ( .D(n70), .CLK(clk), .RSTB(n345), .Q(result[10])
         );
  DFFARX1 \result_reg[9]  ( .D(n69), .CLK(clk), .RSTB(n344), .Q(result[9]) );
  DFFARX1 \result_reg[30]  ( .D(n90), .CLK(clk), .RSTB(n355), .Q(result[30])
         );
  DFFARX1 \result_reg[29]  ( .D(n89), .CLK(clk), .RSTB(n354), .Q(result[29])
         );
  DFFARX1 \result_reg[28]  ( .D(n88), .CLK(clk), .RSTB(n354), .Q(result[28])
         );
  DFFARX1 \result_reg[27]  ( .D(n87), .CLK(clk), .RSTB(n353), .Q(result[27])
         );
  DFFARX1 \result_reg[26]  ( .D(n86), .CLK(clk), .RSTB(n353), .Q(result[26])
         );
  DFFARX1 \result_reg[25]  ( .D(n85), .CLK(clk), .RSTB(n352), .Q(result[25])
         );
  DFFARX1 \result_reg[24]  ( .D(n84), .CLK(clk), .RSTB(n352), .Q(result[24])
         );
  DFFARX1 \result_reg[23]  ( .D(n83), .CLK(clk), .RSTB(n351), .Q(result[23])
         );
  DFFARX1 \result_reg[22]  ( .D(n82), .CLK(clk), .RSTB(n351), .Q(result[22])
         );
  DFFARX1 \result_reg[21]  ( .D(n81), .CLK(clk), .RSTB(n350), .Q(result[21])
         );
  DFFARX1 \result_reg[6]  ( .D(n95), .CLK(clk), .RSTB(n357), .Q(result[6]) );
  DFFARX1 \result_reg[5]  ( .D(n94), .CLK(clk), .RSTB(n357), .Q(result[5]) );
  DFFARX1 \result_reg[4]  ( .D(n93), .CLK(clk), .RSTB(n356), .Q(result[4]) );
  DFFARX1 \result_reg[3]  ( .D(n92), .CLK(clk), .RSTB(n356), .Q(result[3]) );
  DFFARX1 \result_reg[2]  ( .D(n91), .CLK(clk), .RSTB(n355), .Q(result[2]) );
  DFFARX1 \result_reg[0]  ( .D(n99), .CLK(clk), .RSTB(n359), .Q(result[0]) );
  DFFARX1 \reg_a_reg[26]  ( .D(N85), .CLK(clk), .RSTB(n353), .Q(reg_a[26]), 
        .QN(n534) );
  DFFARX1 \reg_b_reg[23]  ( .D(N115), .CLK(clk), .RSTB(n351), .Q(reg_b[23]), 
        .QN(n371) );
  DFFARX1 \reg_b_reg[17]  ( .D(N109), .CLK(clk), .RSTB(n348), .Q(reg_b[17]), 
        .QN(n377) );
  DFFARX1 \reg_b_reg[31]  ( .D(N123), .CLK(clk), .RSTB(n358), .Q(reg_b[31]), 
        .QN(n586) );
  DFFARX1 \reg_b_reg[28]  ( .D(N120), .CLK(clk), .RSTB(n354), .Q(reg_b[28]) );
  DFFARX1 \reg_b_reg[27]  ( .D(N119), .CLK(clk), .RSTB(n353), .Q(reg_b[27]) );
  DFFARX1 \reg_b_reg[13]  ( .D(N105), .CLK(clk), .RSTB(n346), .Q(reg_b[13]), 
        .QN(n383) );
  DFFARX1 \reg_b_reg[26]  ( .D(N118), .CLK(clk), .RSTB(n353), .Q(reg_b[26]), 
        .QN(n370) );
  DFFARX1 \reg_b_reg[14]  ( .D(N106), .CLK(clk), .RSTB(n347), .Q(reg_b[14]), 
        .QN(n380) );
  DFFARX1 \reg_b_reg[11]  ( .D(N103), .CLK(clk), .RSTB(n345), .Q(reg_b[11]), 
        .QN(n384) );
  DFFARX1 \reg_b_reg[20]  ( .D(N112), .CLK(clk), .RSTB(n350), .Q(reg_b[20]), 
        .QN(n374) );
  DFFARX1 \reg_b_reg[3]  ( .D(N95), .CLK(clk), .RSTB(n356), .Q(reg_b[3]) );
  DFFARX1 \reg_a_reg[30]  ( .D(N89), .CLK(clk), .RSTB(n355), .Q(reg_a[30]) );
  DFFARX1 \reg_a_reg[29]  ( .D(N88), .CLK(clk), .RSTB(n354), .Q(reg_a[29]) );
  DFFARX1 \reg_a_reg[11]  ( .D(N70), .CLK(clk), .RSTB(n345), .Q(reg_a[11]) );
  DFFARX1 \reg_a_reg[9]  ( .D(N68), .CLK(clk), .RSTB(n344), .Q(reg_a[9]) );
  DFFARX1 \reg_a_reg[10]  ( .D(N69), .CLK(clk), .RSTB(n345), .Q(reg_a[10]) );
  DFFARX1 \reg_a_reg[27]  ( .D(N86), .CLK(clk), .RSTB(n353), .Q(reg_a[27]), 
        .QN(n423) );
  DFFARX1 \reg_a_reg[23]  ( .D(N82), .CLK(clk), .RSTB(n351), .Q(reg_a[23]) );
  DFFARX1 \reg_a_reg[22]  ( .D(N81), .CLK(clk), .RSTB(n351), .Q(reg_a[22]) );
  DFFARX1 \reg_a_reg[14]  ( .D(N73), .CLK(clk), .RSTB(n347), .Q(reg_a[14]) );
  DFFARX1 \reg_a_reg[25]  ( .D(N84), .CLK(clk), .RSTB(n352), .Q(reg_a[25]) );
  DFFARX1 \reg_b_reg[5]  ( .D(N97), .CLK(clk), .RSTB(n357), .Q(n119), .QN(n240) );
  DFFARX1 \reg_a_reg[6]  ( .D(N65), .CLK(clk), .RSTB(n357), .QN(n157) );
  DFFARX1 \reg_a_reg[1]  ( .D(N60), .CLK(clk), .RSTB(n359), .QN(n163) );
  DFFARX1 \reg_a_reg[17]  ( .D(N76), .CLK(clk), .RSTB(n348), .Q(reg_a[17]) );
  DFFARX2 \reg_a_reg[7]  ( .D(N66), .CLK(clk), .RSTB(n358), .QN(n150) );
  OR2X2 U166 ( .IN1(reg_a[9]), .IN2(n228), .Q(n450) );
  OR2X1 U167 ( .IN1(n398), .IN2(n575), .Q(n440) );
  NAND2X2 U168 ( .IN1(n125), .IN2(n126), .QN(n575) );
  INVX4 U169 ( .IN(n200), .QN(n608) );
  INVX2 U170 ( .IN(reg_a[17]), .QN(n102) );
  INVX4 U171 ( .IN(n102), .QN(n103) );
  INVX8 U172 ( .IN(n444), .QN(n104) );
  INVX16 U173 ( .IN(n104), .QN(n105) );
  INVX4 U174 ( .IN(n208), .QN(n153) );
  INVX8 U175 ( .IN(n191), .QN(n146) );
  NOR2X4 U176 ( .IN1(n269), .IN2(n600), .QN(n191) );
  NOR2X0 U177 ( .IN1(n387), .IN2(n172), .QN(n131) );
  INVX0 U178 ( .IN(n396), .QN(n387) );
  NOR2X0 U179 ( .IN1(n525), .IN2(n110), .QN(n415) );
  INVX0 U180 ( .IN(n509), .QN(n372) );
  INVX0 U181 ( .IN(n209), .QN(n154) );
  NAND2X2 U182 ( .IN1(n152), .IN2(n241), .QN(n570) );
  OR2X1 U183 ( .IN1(n232), .IN2(n240), .Q(n396) );
  OR2X1 U184 ( .IN1(reg_a[14]), .IN2(n380), .Q(n382) );
  OR2X1 U185 ( .IN1(reg_a[11]), .IN2(n384), .Q(n386) );
  INVX0 U186 ( .IN(n386), .QN(n405) );
  OR2X1 U187 ( .IN1(n122), .IN2(n161), .Q(n138) );
  NAND2X0 U188 ( .IN1(n218), .IN2(reg_b[24]), .QN(n518) );
  INVX0 U189 ( .IN(n497), .QN(n272) );
  NAND2X0 U190 ( .IN1(n221), .IN2(reg_b[21]), .QN(n504) );
  NAND2X1 U191 ( .IN1(n164), .IN2(n440), .QN(n399) );
  AND2X1 U192 ( .IN1(n131), .IN2(n164), .Q(n166) );
  NAND2X2 U193 ( .IN1(n451), .IN2(n108), .QN(n403) );
  OR2X1 U194 ( .IN1(n211), .IN2(reg_b[28]), .Q(n426) );
  INVX0 U195 ( .IN(n514), .QN(n144) );
  OR2X1 U196 ( .IN1(n599), .IN2(n436), .Q(n249) );
  OR2X1 U197 ( .IN1(reg_a[20]), .IN2(n374), .Q(n376) );
  AO22X1 U198 ( .IN1(n375), .IN2(n376), .IN3(reg_a[20]), .IN4(n374), .Q(n501)
         );
  INVX0 U199 ( .IN(n496), .QN(n375) );
  NAND2X0 U200 ( .IN1(n224), .IN2(reg_b[12]), .QN(n464) );
  NAND2X0 U201 ( .IN1(n219), .IN2(reg_b[18]), .QN(n491) );
  NAND2X0 U202 ( .IN1(n212), .IN2(n100), .QN(n436) );
  OR2X1 U203 ( .IN1(n599), .IN2(n436), .Q(n434) );
  OR2X1 U204 ( .IN1(n395), .IN2(n442), .Q(n447) );
  OR2X1 U205 ( .IN1(n599), .IN2(n436), .Q(n200) );
  NOR4X0 U206 ( .IN1(n65), .IN2(n66), .IN3(n63), .IN4(n64), .QN(n186) );
  NOR4X0 U207 ( .IN1(n61), .IN2(n62), .IN3(n59), .IN4(n60), .QN(n187) );
  NAND2X1 U208 ( .IN1(n209), .IN2(n155), .QN(n441) );
  NAND2X2 U209 ( .IN1(n139), .IN2(n578), .QN(n442) );
  NAND2X0 U210 ( .IN1(n150), .IN2(n112), .QN(n139) );
  INVX2 U211 ( .IN(n129), .QN(n151) );
  OA21X1 U212 ( .IN1(n114), .IN2(n554), .IN3(n553), .Q(n195) );
  INVX0 U213 ( .IN(n414), .QN(n515) );
  NAND2X0 U214 ( .IN1(n213), .IN2(reg_a[15]), .QN(n479) );
  NAND2X0 U215 ( .IN1(n214), .IN2(reg_a[18]), .QN(n492) );
  NOR2X0 U216 ( .IN1(n170), .IN2(n118), .QN(n169) );
  NAND2X2 U217 ( .IN1(n210), .IN2(n153), .QN(n563) );
  NAND2X0 U218 ( .IN1(n215), .IN2(reg_a[12]), .QN(n465) );
  NBUFFX2 U219 ( .IN(n604), .Q(n284) );
  INVX0 U220 ( .IN(n134), .QN(n498) );
  NAND2X0 U221 ( .IN1(n216), .IN2(reg_a[19]), .QN(n496) );
  OAI21X1 U222 ( .IN1(reg_a[19]), .IN2(n216), .IN3(n491), .QN(n497) );
  INVX4 U223 ( .IN(n146), .QN(n148) );
  INVX4 U224 ( .IN(n146), .QN(n147) );
  INVX4 U225 ( .IN(n146), .QN(n149) );
  XOR3X1 U226 ( .IN1(reg_b[17]), .IN2(n103), .IN3(n485), .Q(n487) );
  XOR3X1 U227 ( .IN1(n237), .IN2(n113), .IN3(n194), .Q(n577) );
  XOR3X1 U228 ( .IN1(reg_b[27]), .IN2(reg_a[27]), .IN3(n539), .Q(n541) );
  NAND2X0 U229 ( .IN1(n538), .IN2(n537), .QN(N85) );
  NOR2X0 U230 ( .IN1(n536), .IN2(n535), .QN(n537) );
  NAND2X0 U231 ( .IN1(n598), .IN2(n597), .QN(N60) );
  NOR2X0 U232 ( .IN1(n596), .IN2(n595), .QN(n597) );
  XOR3X1 U233 ( .IN1(n154), .IN2(n155), .IN3(n581), .Q(n583) );
  INVX0 U234 ( .IN(n165), .QN(n542) );
  AND2X1 U235 ( .IN1(n207), .IN2(n599), .Q(gcd_ns[1]) );
  XOR3X1 U236 ( .IN1(n232), .IN2(n119), .IN3(n572), .Q(n574) );
  NAND2X4 U237 ( .IN1(n159), .IN2(reg_b[1]), .QN(n160) );
  AND2X1 U238 ( .IN1(n558), .IN2(n559), .Q(n201) );
  NAND2X0 U239 ( .IN1(n559), .IN2(n563), .QN(n388) );
  NAND2X1 U240 ( .IN1(n243), .IN2(n242), .QN(n559) );
  INVX8 U241 ( .IN(n600), .QN(n277) );
  NOR2X0 U242 ( .IN1(reg_a[30]), .IN2(n223), .QN(n107) );
  AOI22X1 U243 ( .IN1(n402), .IN2(n401), .IN3(n151), .IN4(n130), .QN(n108) );
  INVX2 U244 ( .IN(n105), .QN(n145) );
  INVX2 U245 ( .IN(n277), .QN(n276) );
  NOR2X0 U246 ( .IN1(reg_a[26]), .IN2(n370), .QN(n110) );
  AND2X1 U247 ( .IN1(n196), .IN2(n373), .Q(n111) );
  AND2X1 U248 ( .IN1(n426), .IN2(n425), .Q(n114) );
  OR2X1 U249 ( .IN1(n471), .IN2(n407), .Q(n115) );
  AND2X1 U250 ( .IN1(n272), .IN2(n376), .Q(n116) );
  OR2X1 U251 ( .IN1(reg_b[27]), .IN2(n423), .Q(n117) );
  OR2X1 U252 ( .IN1(n484), .IN2(n409), .Q(n118) );
  NAND2X0 U253 ( .IN1(n186), .IN2(n187), .QN(n6) );
  OR2X1 U254 ( .IN1(n461), .IN2(n406), .Q(n120) );
  AND2X1 U255 ( .IN1(n246), .IN2(n505), .Q(n121) );
  OR2X1 U256 ( .IN1(n475), .IN2(n408), .Q(n122) );
  INVX2 U257 ( .IN(n157), .QN(n237) );
  AOI22X1 U258 ( .IN1(n168), .IN2(reg_b[30]), .IN3(n234), .IN4(reg_a[30]), 
        .QN(n123) );
  INVX2 U259 ( .IN(n150), .QN(n155) );
  INVX2 U260 ( .IN(n163), .QN(n242) );
  INVX0 U261 ( .IN(n242), .QN(n159) );
  NOR2X0 U262 ( .IN1(n404), .IN2(n403), .QN(n124) );
  OR2X2 U263 ( .IN1(n488), .IN2(n410), .Q(n161) );
  INVX8 U264 ( .IN(n127), .QN(n599) );
  NAND2X1 U265 ( .IN1(n397), .IN2(n396), .QN(n125) );
  NAND2X0 U266 ( .IN1(n232), .IN2(n240), .QN(n126) );
  NAND2X4 U267 ( .IN1(n431), .IN2(n432), .QN(n127) );
  OR2X1 U268 ( .IN1(n436), .IN2(n433), .Q(n128) );
  NAND2X2 U269 ( .IN1(n128), .IN2(n435), .QN(n235) );
  INVX0 U270 ( .IN(n570), .QN(n397) );
  INVX2 U271 ( .IN(n156), .QN(n232) );
  NAND2X2 U272 ( .IN1(n431), .IN2(n432), .QN(n433) );
  OR2X1 U273 ( .IN1(n607), .IN2(n231), .Q(n435) );
  NOR2X0 U274 ( .IN1(n199), .IN2(n122), .QN(n170) );
  NOR2X0 U275 ( .IN1(n241), .IN2(n152), .QN(n172) );
  NAND2X0 U276 ( .IN1(n529), .IN2(n528), .QN(n530) );
  NAND2X0 U277 ( .IN1(n288), .IN2(n557), .QN(n132) );
  NAND2X0 U278 ( .IN1(a_in[30]), .IN2(n280), .QN(n133) );
  NAND3X0 U279 ( .IN1(n132), .IN2(n133), .IN3(n123), .QN(N89) );
  DELLN1X2 U280 ( .IN(n411), .Q(n134) );
  NBUFFX16 U281 ( .IN(n606), .Q(n288) );
  NBUFFX16 U282 ( .IN(n604), .Q(n280) );
  NOR2X4 U283 ( .IN1(n199), .IN2(n138), .QN(n135) );
  NOR2X4 U284 ( .IN1(n135), .IN2(n136), .QN(n411) );
  AND2X1 U285 ( .IN1(n137), .IN2(n118), .Q(n136) );
  INVX0 U286 ( .IN(n161), .QN(n137) );
  OR4X4 U287 ( .IN1(reg_b[31]), .IN2(reg_b[3]), .IN3(n109), .IN4(n119), .Q(n60) );
  NAND2X4 U288 ( .IN1(n392), .IN2(n562), .QN(n394) );
  NOR2X4 U289 ( .IN1(n391), .IN2(n390), .QN(n392) );
  NOR2X4 U290 ( .IN1(n389), .IN2(n388), .QN(n391) );
  OR2X2 U291 ( .IN1(n127), .IN2(n436), .Q(n140) );
  NAND2X4 U292 ( .IN1(n140), .IN2(n435), .QN(n600) );
  INVX4 U293 ( .IN(n277), .QN(n275) );
  NOR2X4 U294 ( .IN1(n599), .IN2(n436), .QN(n248) );
  NAND2X4 U295 ( .IN1(n600), .IN2(n145), .QN(n141) );
  INVX2 U296 ( .IN(n401), .QN(n395) );
  NOR2X2 U297 ( .IN1(n534), .IN2(n239), .QN(n536) );
  INVX8 U298 ( .IN(n591), .QN(n606) );
  NAND2X4 U299 ( .IN1(n600), .IN2(n105), .QN(n591) );
  NAND2X4 U300 ( .IN1(n143), .IN2(n142), .QN(n429) );
  OR2X1 U301 ( .IN1(n545), .IN2(n427), .Q(n142) );
  NOR2X4 U302 ( .IN1(n428), .IN2(n107), .QN(n143) );
  NAND2X4 U303 ( .IN1(n416), .IN2(n417), .QN(n418) );
  NAND2X2 U304 ( .IN1(n415), .IN2(n527), .QN(n416) );
  NAND3X0 U305 ( .IN1(n414), .IN2(n144), .IN3(n519), .QN(n527) );
  NAND2X4 U306 ( .IN1(n166), .IN2(n438), .QN(n400) );
  NAND2X2 U307 ( .IN1(n105), .IN2(n277), .QN(n590) );
  OR2X2 U308 ( .IN1(n151), .IN2(n130), .Q(n401) );
  OR4X2 U309 ( .IN1(n113), .IN2(n154), .IN3(n106), .IN4(reg_b[9]), .Q(n59) );
  OR2X2 U310 ( .IN1(n113), .IN2(n157), .Q(n579) );
  IBUFFX16 U311 ( .IN(n578), .QN(n580) );
  NAND2X4 U312 ( .IN1(n399), .IN2(n400), .QN(n404) );
  NAND2X4 U313 ( .IN1(n197), .IN2(n111), .QN(n414) );
  OR2X2 U314 ( .IN1(n237), .IN2(n236), .Q(n578) );
  NOR2X4 U315 ( .IN1(n105), .IN2(n235), .QN(n158) );
  NAND2X4 U316 ( .IN1(n160), .IN2(n601), .QN(n558) );
  INVX4 U317 ( .IN(n558), .QN(n389) );
  OR2X1 U318 ( .IN1(n437), .IN2(n207), .Q(n162) );
  NOR2X4 U319 ( .IN1(n248), .IN2(n162), .QN(n444) );
  INVX0 U320 ( .IN(n435), .QN(n437) );
  NOR2X0 U321 ( .IN1(n6), .IN2(n436), .QN(n207) );
  NAND2X4 U322 ( .IN1(n411), .IN2(n116), .QN(n247) );
  NAND2X4 U323 ( .IN1(n247), .IN2(n121), .QN(n197) );
  NOR2X4 U324 ( .IN1(n395), .IN2(n442), .QN(n164) );
  NAND2X4 U325 ( .IN1(n422), .IN2(n117), .QN(n165) );
  INVX0 U326 ( .IN(n501), .QN(n246) );
  NAND2X0 U327 ( .IN1(n227), .IN2(reg_a[21]), .QN(n505) );
  NOR2X4 U328 ( .IN1(n171), .IN2(n115), .QN(n199) );
  INVX0 U329 ( .IN(n382), .QN(n407) );
  OR2X1 U330 ( .IN1(reg_a[23]), .IN2(n371), .Q(n373) );
  NOR2X0 U331 ( .IN1(n529), .IN2(n110), .QN(n419) );
  NAND2X2 U332 ( .IN1(n225), .IN2(reg_a[10]), .QN(n455) );
  INVX0 U333 ( .IN(n249), .QN(n268) );
  NOR2X4 U334 ( .IN1(n404), .IN2(n403), .QN(n457) );
  OA21X1 U335 ( .IN1(n520), .IN2(n203), .IN3(n519), .Q(n521) );
  OA21X1 U336 ( .IN1(n271), .IN2(n510), .IN3(n509), .Q(n511) );
  NAND2X0 U337 ( .IN1(n228), .IN2(reg_a[9]), .QN(n451) );
  INVX2 U338 ( .IN(n483), .QN(n378) );
  OAI21X1 U339 ( .IN1(reg_a[22]), .IN2(n229), .IN3(n504), .QN(n510) );
  NOR2X4 U340 ( .IN1(n198), .IN2(n120), .QN(n171) );
  IBUFFX2 U341 ( .IN(n379), .QN(n409) );
  NOR2X4 U342 ( .IN1(n105), .IN2(n235), .QN(n167) );
  NOR2X4 U343 ( .IN1(n105), .IN2(n235), .QN(n168) );
  NBUFFX2 U344 ( .IN(n604), .Q(n279) );
  INVX2 U345 ( .IN(n249), .QN(n269) );
  INVX0 U346 ( .IN(n105), .QN(n192) );
  INVX0 U347 ( .IN(n510), .QN(n196) );
  NOR2X0 U348 ( .IN1(n274), .IN2(n501), .QN(n173) );
  NOR2X2 U349 ( .IN1(n456), .IN2(n405), .QN(n188) );
  INVX2 U350 ( .IN(n188), .QN(n189) );
  AND2X1 U351 ( .IN1(n183), .IN2(reg_b[3]), .Q(n390) );
  NAND2X0 U352 ( .IN1(reg_b[31]), .IN2(n174), .QN(n432) );
  XOR3X1 U353 ( .IN1(n225), .IN2(reg_a[10]), .IN3(n175), .Q(n454) );
  OAI21X1 U354 ( .IN1(n452), .IN2(n202), .IN3(n451), .QN(n175) );
  XOR3X1 U355 ( .IN1(n176), .IN2(reg_a[16]), .IN3(n177), .Q(n482) );
  OAI21X1 U356 ( .IN1(n480), .IN2(n206), .IN3(n479), .QN(n177) );
  XOR3X1 U357 ( .IN1(reg_b[19]), .IN2(n178), .IN3(n179), .Q(n495) );
  OAI21X1 U358 ( .IN1(n493), .IN2(n204), .IN3(n492), .QN(n179) );
  XOR3X1 U359 ( .IN1(reg_b[20]), .IN2(n180), .IN3(n181), .Q(n500) );
  OAI21X1 U360 ( .IN1(n498), .IN2(n497), .IN3(n496), .QN(n181) );
  XOR3X1 U361 ( .IN1(n229), .IN2(reg_a[22]), .IN3(n182), .Q(n508) );
  OAI21X1 U362 ( .IN1(n506), .IN2(n173), .IN3(n505), .QN(n182) );
  OR2X1 U363 ( .IN1(n183), .IN2(reg_b[3]), .Q(n393) );
  NAND2X4 U364 ( .IN1(n220), .IN2(reg_b[15]), .QN(n478) );
  OR2X1 U365 ( .IN1(reg_b[13]), .IN2(n184), .Q(n470) );
  OAI21X1 U366 ( .IN1(reg_a[10]), .IN2(n225), .IN3(n450), .QN(n456) );
  OR2X1 U367 ( .IN1(reg_b[16]), .IN2(n185), .Q(n483) );
  NAND2X0 U368 ( .IN1(reg_b[28]), .IN2(n211), .QN(n424) );
  NOR2X4 U369 ( .IN1(n457), .IN2(n189), .QN(n198) );
  NBUFFX2 U370 ( .IN(n606), .Q(n287) );
  NBUFFX2 U371 ( .IN(n606), .Q(n289) );
  NBUFFX2 U372 ( .IN(n606), .Q(n286) );
  NBUFFX2 U373 ( .IN(n604), .Q(n278) );
  NBUFFX2 U374 ( .IN(n604), .Q(n283) );
  NBUFFX2 U375 ( .IN(n604), .Q(n282) );
  NBUFFX2 U376 ( .IN(n604), .Q(n281) );
  NBUFFX2 U377 ( .IN(n606), .Q(n293) );
  NBUFFX2 U378 ( .IN(n604), .Q(n285) );
  INVX0 U379 ( .IN(n327), .QN(n317) );
  INVX0 U380 ( .IN(n326), .QN(n319) );
  INVX0 U381 ( .IN(n327), .QN(n318) );
  INVX0 U382 ( .IN(n326), .QN(n320) );
  NBUFFX2 U383 ( .IN(n606), .Q(n292) );
  NBUFFX2 U384 ( .IN(n606), .Q(n291) );
  NBUFFX2 U385 ( .IN(n606), .Q(n290) );
  INVX0 U386 ( .IN(n325), .QN(n322) );
  INVX0 U387 ( .IN(n324), .QN(n323) );
  INVX0 U388 ( .IN(n325), .QN(n321) );
  INVX0 U389 ( .IN(n303), .QN(n327) );
  INVX0 U390 ( .IN(n303), .QN(n326) );
  INVX0 U391 ( .IN(n6), .QN(n328) );
  INVX0 U392 ( .IN(n310), .QN(n329) );
  INVX0 U393 ( .IN(n304), .QN(n330) );
  INVX0 U394 ( .IN(n305), .QN(n332) );
  INVX0 U395 ( .IN(n305), .QN(n333) );
  INVX0 U396 ( .IN(n306), .QN(n334) );
  INVX0 U397 ( .IN(n306), .QN(n335) );
  INVX0 U398 ( .IN(n307), .QN(n336) );
  INVX0 U399 ( .IN(n307), .QN(n337) );
  INVX0 U400 ( .IN(n308), .QN(n338) );
  INVX0 U401 ( .IN(n308), .QN(n339) );
  INVX0 U402 ( .IN(n309), .QN(n340) );
  INVX0 U403 ( .IN(n304), .QN(n331) );
  INVX0 U404 ( .IN(n310), .QN(n343) );
  INVX0 U405 ( .IN(n309), .QN(n341) );
  INVX0 U406 ( .IN(n310), .QN(n342) );
  NOR2X0 U407 ( .IN1(n193), .IN2(n440), .QN(n190) );
  INVX0 U408 ( .IN(n579), .QN(n398) );
  OR2X1 U409 ( .IN1(n387), .IN2(n172), .Q(n439) );
  NAND2X4 U410 ( .IN1(n275), .IN2(n192), .QN(n239) );
  INVX0 U411 ( .IN(n302), .QN(n324) );
  INVX0 U412 ( .IN(n315), .QN(n303) );
  INVX0 U413 ( .IN(n314), .QN(n304) );
  INVX0 U414 ( .IN(n314), .QN(n305) );
  INVX0 U415 ( .IN(n302), .QN(n325) );
  INVX0 U416 ( .IN(n313), .QN(n306) );
  INVX0 U417 ( .IN(n313), .QN(n307) );
  INVX0 U418 ( .IN(n312), .QN(n308) );
  INVX0 U419 ( .IN(n312), .QN(n309) );
  INVX0 U420 ( .IN(n311), .QN(n310) );
  OR2X1 U421 ( .IN1(n552), .IN2(n546), .Q(n427) );
  NOR2X0 U422 ( .IN1(n571), .IN2(n439), .QN(n193) );
  NOR2X0 U423 ( .IN1(n193), .IN2(n575), .QN(n194) );
  INVX0 U424 ( .IN(n434), .QN(n266) );
  INVX0 U425 ( .IN(n434), .QN(n267) );
  OR2X1 U426 ( .IN1(n546), .IN2(n554), .Q(n549) );
  OR2X1 U427 ( .IN1(n552), .IN2(n107), .Q(n556) );
  INVX0 U428 ( .IN(n492), .QN(n410) );
  NOR2X0 U429 ( .IN1(n594), .IN2(n593), .QN(n598) );
  NOR2X0 U430 ( .IN1(n590), .IN2(n589), .QN(n594) );
  INVX0 U431 ( .IN(n479), .QN(n408) );
  INVX0 U432 ( .IN(n465), .QN(n406) );
  NOR2X0 U433 ( .IN1(n533), .IN2(n532), .QN(n538) );
  NOR2X0 U434 ( .IN1(n590), .IN2(n524), .QN(n533) );
  INVX0 U435 ( .IN(n505), .QN(n413) );
  INVX0 U436 ( .IN(n6), .QN(n315) );
  INVX0 U437 ( .IN(n6), .QN(n314) );
  INVX0 U438 ( .IN(n6), .QN(n313) );
  INVX0 U439 ( .IN(n6), .QN(n312) );
  INVX0 U440 ( .IN(n6), .QN(n311) );
  INVX0 U441 ( .IN(n316), .QN(n302) );
  INVX0 U442 ( .IN(n6), .QN(n316) );
  INVX0 U443 ( .IN(n438), .QN(n571) );
  OR3X1 U444 ( .IN1(n231), .IN2(n609), .IN3(n262), .Q(gcd_ns[0]) );
  AND2X1 U445 ( .IN1(n607), .IN2(n308), .Q(n609) );
  OA21X1 U446 ( .IN1(n190), .IN2(n447), .IN3(n108), .Q(n202) );
  INVX0 U447 ( .IN(n436), .QN(n607) );
  INVX0 U448 ( .IN(n525), .QN(n526) );
  INVX0 U449 ( .IN(n545), .QN(n554) );
  INVX0 U450 ( .IN(n553), .QN(n546) );
  INVX0 U451 ( .IN(n584), .QN(n552) );
  NOR2X0 U452 ( .IN1(n515), .IN2(n514), .QN(n203) );
  NOR2X0 U453 ( .IN1(n169), .IN2(n488), .QN(n204) );
  NOR2X0 U454 ( .IN1(n198), .IN2(n461), .QN(n205) );
  NOR2X0 U455 ( .IN1(n199), .IN2(n475), .QN(n206) );
  INVX0 U456 ( .IN(n376), .QN(n412) );
  INVX0 U457 ( .IN(n562), .QN(n564) );
  INVX0 U458 ( .IN(n450), .QN(n452) );
  INVX0 U459 ( .IN(n478), .QN(n480) );
  INVX0 U460 ( .IN(n491), .QN(n493) );
  INVX0 U461 ( .IN(n504), .QN(n506) );
  INVX0 U462 ( .IN(n518), .QN(n520) );
  INVX0 U463 ( .IN(n464), .QN(n466) );
  NBUFFX2 U464 ( .IN(n362), .Q(n357) );
  NBUFFX2 U465 ( .IN(n361), .Q(n359) );
  NBUFFX2 U466 ( .IN(n363), .Q(n356) );
  NBUFFX2 U467 ( .IN(n368), .Q(n345) );
  NBUFFX2 U468 ( .IN(n368), .Q(n346) );
  NBUFFX2 U469 ( .IN(n367), .Q(n347) );
  NBUFFX2 U470 ( .IN(n367), .Q(n348) );
  NBUFFX2 U471 ( .IN(n366), .Q(n349) );
  NBUFFX2 U472 ( .IN(n366), .Q(n350) );
  NBUFFX2 U473 ( .IN(n365), .Q(n351) );
  NBUFFX2 U474 ( .IN(n365), .Q(n352) );
  NBUFFX2 U475 ( .IN(n364), .Q(n353) );
  NBUFFX2 U476 ( .IN(n364), .Q(n354) );
  NBUFFX2 U477 ( .IN(n363), .Q(n355) );
  NBUFFX2 U478 ( .IN(n362), .Q(n358) );
  NBUFFX2 U479 ( .IN(n361), .Q(n360) );
  INVX0 U480 ( .IN(n441), .QN(n402) );
  AO222X1 U481 ( .IN1(n268), .IN2(reg_a[31]), .IN3(b_in[31]), .IN4(n148), 
        .IN5(reg_b[31]), .IN6(n276), .Q(N123) );
  AO222X1 U482 ( .IN1(n252), .IN2(reg_a[20]), .IN3(b_in[20]), .IN4(n149), 
        .IN5(reg_b[20]), .IN6(n276), .Q(N112) );
  AO222X1 U483 ( .IN1(n250), .IN2(reg_a[22]), .IN3(b_in[22]), .IN4(n148), 
        .IN5(reg_b[22]), .IN6(n275), .Q(N114) );
  AO222X1 U484 ( .IN1(n267), .IN2(reg_a[23]), .IN3(b_in[23]), .IN4(n149), 
        .IN5(reg_b[23]), .IN6(n276), .Q(N115) );
  AO222X1 U485 ( .IN1(n269), .IN2(reg_a[10]), .IN3(b_in[10]), .IN4(n148), 
        .IN5(reg_b[10]), .IN6(n276), .Q(N102) );
  AO222X1 U486 ( .IN1(n260), .IN2(reg_a[11]), .IN3(b_in[11]), .IN4(n148), 
        .IN5(reg_b[11]), .IN6(n275), .Q(N103) );
  AO222X1 U487 ( .IN1(n255), .IN2(reg_a[14]), .IN3(b_in[14]), .IN4(n148), 
        .IN5(reg_b[14]), .IN6(n275), .Q(N106) );
  AO222X1 U488 ( .IN1(n268), .IN2(reg_a[15]), .IN3(b_in[15]), .IN4(n148), 
        .IN5(reg_b[15]), .IN6(n275), .Q(N107) );
  AO222X1 U489 ( .IN1(n266), .IN2(reg_a[16]), .IN3(b_in[16]), .IN4(n147), 
        .IN5(reg_b[16]), .IN6(n276), .Q(N108) );
  AO222X1 U490 ( .IN1(n269), .IN2(n103), .IN3(b_in[17]), .IN4(n148), .IN5(
        reg_b[17]), .IN6(n276), .Q(N109) );
  AO222X1 U491 ( .IN1(n253), .IN2(reg_a[25]), .IN3(b_in[25]), .IN4(n148), 
        .IN5(reg_b[25]), .IN6(n275), .Q(N117) );
  AO222X1 U492 ( .IN1(n259), .IN2(reg_a[27]), .IN3(b_in[27]), .IN4(n149), 
        .IN5(reg_b[27]), .IN6(n275), .Q(N119) );
  AO222X1 U493 ( .IN1(n257), .IN2(reg_a[29]), .IN3(b_in[29]), .IN4(n147), 
        .IN5(reg_b[29]), .IN6(n276), .Q(N121) );
  AO222X1 U494 ( .IN1(n252), .IN2(reg_a[3]), .IN3(b_in[3]), .IN4(n147), .IN5(
        reg_b[3]), .IN6(n275), .Q(N95) );
  NAND2X0 U495 ( .IN1(n208), .IN2(reg_b[2]), .QN(n562) );
  AND3X1 U496 ( .IN1(reg_a[31]), .IN2(n586), .IN3(n585), .Q(n588) );
  OAI21X1 U497 ( .IN1(n107), .IN2(n195), .IN3(n584), .QN(n585) );
  MUX21X1 U498 ( .IN1(n549), .IN2(n548), .S(n114), .Q(n551) );
  XOR2X1 U499 ( .IN1(n222), .IN2(reg_a[29]), .Q(n548) );
  XOR3X1 U500 ( .IN1(reg_b[3]), .IN2(reg_a[3]), .IN3(n565), .Q(n567) );
  OA21X1 U501 ( .IN1(n564), .IN2(n201), .IN3(n563), .Q(n565) );
  XOR3X1 U502 ( .IN1(reg_b[25]), .IN2(reg_a[25]), .IN3(n521), .Q(n523) );
  XOR3X1 U503 ( .IN1(n153), .IN2(reg_b[2]), .IN3(n201), .Q(n561) );
  XOR3X1 U504 ( .IN1(reg_b[14]), .IN2(reg_a[14]), .IN3(n472), .Q(n474) );
  XOR3X1 U505 ( .IN1(reg_b[23]), .IN2(reg_a[23]), .IN3(n511), .Q(n513) );
  XOR3X1 U506 ( .IN1(n106), .IN2(n151), .IN3(n443), .Q(n446) );
  AND2X1 U507 ( .IN1(reg_b[1]), .IN2(n168), .Q(n595) );
  AND2X1 U508 ( .IN1(reg_b[26]), .IN2(n167), .Q(n535) );
  XOR3X1 U509 ( .IN1(reg_b[28]), .IN2(reg_a[28]), .IN3(n542), .Q(n544) );
  MUX21X1 U510 ( .IN1(n556), .IN2(n555), .S(n195), .Q(n557) );
  XOR2X1 U511 ( .IN1(n223), .IN2(reg_a[30]), .Q(n555) );
  XOR3X1 U512 ( .IN1(reg_a[12]), .IN2(reg_b[12]), .IN3(n205), .Q(n463) );
  XOR3X1 U513 ( .IN1(reg_a[15]), .IN2(reg_b[15]), .IN3(n206), .Q(n477) );
  XOR3X1 U514 ( .IN1(reg_a[9]), .IN2(reg_b[9]), .IN3(n202), .Q(n449) );
  XOR3X1 U515 ( .IN1(reg_a[18]), .IN2(reg_b[18]), .IN3(n204), .Q(n490) );
  XOR3X1 U516 ( .IN1(reg_a[21]), .IN2(reg_b[21]), .IN3(n173), .Q(n503) );
  XOR3X1 U517 ( .IN1(reg_a[24]), .IN2(reg_b[24]), .IN3(n203), .Q(n517) );
  OA21X1 U518 ( .IN1(n466), .IN2(n205), .IN3(n465), .Q(n467) );
  OA21X1 U519 ( .IN1(n580), .IN2(n194), .IN3(n579), .Q(n581) );
  XOR3X1 U520 ( .IN1(reg_b[11]), .IN2(reg_a[11]), .IN3(n458), .Q(n460) );
  OAI21X1 U521 ( .IN1(reg_b[0]), .IN2(n244), .IN3(n601), .QN(n605) );
  INVX4 U522 ( .IN(n238), .QN(n241) );
  NAND2X2 U523 ( .IN1(n394), .IN2(n393), .QN(n438) );
  XOR3X1 U524 ( .IN1(reg_b[26]), .IN2(reg_a[26]), .IN3(n530), .Q(n531) );
  XOR3X1 U525 ( .IN1(n242), .IN2(n601), .IN3(reg_b[1]), .Q(n592) );
  OAI21X1 U526 ( .IN1(reg_a[25]), .IN2(n226), .IN3(n518), .QN(n525) );
  AO22X1 U527 ( .IN1(n372), .IN2(n373), .IN3(reg_a[23]), .IN4(n371), .Q(n514)
         );
  AO22X1 U528 ( .IN1(n381), .IN2(n382), .IN3(reg_a[14]), .IN4(n380), .Q(n475)
         );
  INVX0 U529 ( .IN(n470), .QN(n381) );
  AO22X1 U530 ( .IN1(n385), .IN2(n386), .IN3(reg_a[11]), .IN4(n384), .Q(n461)
         );
  INVX0 U531 ( .IN(n455), .QN(n385) );
  OR4X1 U532 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n63) );
  OR4X1 U533 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n62) );
  OR4X1 U534 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(
        reg_b[16]), .Q(n65) );
  OR2X1 U535 ( .IN1(reg_a[29]), .IN2(n222), .Q(n545) );
  AO22X1 U536 ( .IN1(n151), .IN2(n328), .IN3(result[8]), .IN4(n304), .Q(n68)
         );
  AO22X1 U537 ( .IN1(reg_a[9]), .IN2(n329), .IN3(result[9]), .IN4(n323), .Q(
        n69) );
  AO22X1 U538 ( .IN1(reg_a[10]), .IN2(n329), .IN3(result[10]), .IN4(n323), .Q(
        n70) );
  AO22X1 U539 ( .IN1(reg_a[11]), .IN2(n330), .IN3(result[11]), .IN4(n323), .Q(
        n71) );
  AO22X1 U540 ( .IN1(reg_a[12]), .IN2(n330), .IN3(result[12]), .IN4(n323), .Q(
        n72) );
  AO22X1 U541 ( .IN1(reg_a[14]), .IN2(n331), .IN3(result[14]), .IN4(n322), .Q(
        n74) );
  AO22X1 U542 ( .IN1(reg_a[15]), .IN2(n332), .IN3(result[15]), .IN4(n322), .Q(
        n75) );
  AO22X1 U543 ( .IN1(reg_a[16]), .IN2(n332), .IN3(result[16]), .IN4(n322), .Q(
        n76) );
  AO22X1 U544 ( .IN1(n103), .IN2(n333), .IN3(result[17]), .IN4(n321), .Q(n77)
         );
  AO22X1 U545 ( .IN1(reg_a[18]), .IN2(n333), .IN3(result[18]), .IN4(n321), .Q(
        n78) );
  AO22X1 U546 ( .IN1(reg_a[19]), .IN2(n334), .IN3(result[19]), .IN4(n321), .Q(
        n79) );
  AO22X1 U547 ( .IN1(reg_a[20]), .IN2(n334), .IN3(result[20]), .IN4(n321), .Q(
        n80) );
  AO22X1 U548 ( .IN1(reg_a[21]), .IN2(n335), .IN3(result[21]), .IN4(n320), .Q(
        n81) );
  AO22X1 U549 ( .IN1(reg_a[22]), .IN2(n335), .IN3(result[22]), .IN4(n320), .Q(
        n82) );
  AO22X1 U550 ( .IN1(reg_a[23]), .IN2(n336), .IN3(result[23]), .IN4(n320), .Q(
        n83) );
  AO22X1 U551 ( .IN1(reg_a[24]), .IN2(n336), .IN3(result[24]), .IN4(n319), .Q(
        n84) );
  AO22X1 U552 ( .IN1(reg_a[25]), .IN2(n337), .IN3(result[25]), .IN4(n319), .Q(
        n85) );
  AO22X1 U553 ( .IN1(reg_a[26]), .IN2(n337), .IN3(result[26]), .IN4(n319), .Q(
        n86) );
  AO22X1 U554 ( .IN1(reg_a[27]), .IN2(n338), .IN3(result[27]), .IN4(n319), .Q(
        n87) );
  AO22X1 U555 ( .IN1(reg_a[28]), .IN2(n338), .IN3(result[28]), .IN4(n318), .Q(
        n88) );
  AO22X1 U556 ( .IN1(reg_a[29]), .IN2(n339), .IN3(result[29]), .IN4(n318), .Q(
        n89) );
  AO22X1 U557 ( .IN1(reg_a[30]), .IN2(n339), .IN3(result[30]), .IN4(n318), .Q(
        n90) );
  AO22X1 U558 ( .IN1(n153), .IN2(n340), .IN3(result[2]), .IN4(n318), .Q(n91)
         );
  AO22X1 U559 ( .IN1(reg_a[3]), .IN2(n340), .IN3(result[3]), .IN4(n317), .Q(
        n92) );
  AO22X1 U560 ( .IN1(reg_a[31]), .IN2(n343), .IN3(result[31]), .IN4(n309), .Q(
        n97) );
  AO22X1 U561 ( .IN1(reg_a[0]), .IN2(n329), .IN3(result[0]), .IN4(n320), .Q(
        n99) );
  OR2X2 U562 ( .IN1(n103), .IN2(n377), .Q(n379) );
  NAND2X0 U563 ( .IN1(n217), .IN2(reg_a[24]), .QN(n519) );
  NAND2X0 U564 ( .IN1(n222), .IN2(reg_a[29]), .QN(n553) );
  NAND2X0 U565 ( .IN1(n223), .IN2(reg_a[30]), .QN(n584) );
  NAND2X0 U566 ( .IN1(reg_a[26]), .IN2(n370), .QN(n417) );
  NAND2X0 U567 ( .IN1(reg_a[31]), .IN2(n586), .QN(n430) );
  NAND2X0 U568 ( .IN1(n226), .IN2(reg_a[25]), .QN(n529) );
  NAND2X0 U569 ( .IN1(reg_b[27]), .IN2(n423), .QN(n421) );
  OAI21X1 U570 ( .IN1(reg_a[16]), .IN2(n176), .IN3(n478), .QN(n484) );
  INVX0 U571 ( .IN(a_in[1]), .QN(n589) );
  INVX0 U572 ( .IN(a_in[26]), .QN(n524) );
  NAND2X0 U573 ( .IN1(n229), .IN2(reg_a[22]), .QN(n509) );
  AND2X1 U574 ( .IN1(n230), .IN2(n67), .Q(done) );
  AND3X1 U575 ( .IN1(start), .IN2(n67), .IN3(n100), .Q(n231) );
  AO22X1 U576 ( .IN1(n378), .IN2(n379), .IN3(n103), .IN4(n377), .Q(n488) );
  NBUFFX2 U577 ( .IN(n369), .Q(n344) );
  NBUFFX2 U578 ( .IN(reset_n), .Q(n369) );
  NBUFFX2 U579 ( .IN(reset_n), .Q(n368) );
  NBUFFX2 U580 ( .IN(reset_n), .Q(n367) );
  NBUFFX2 U581 ( .IN(reset_n), .Q(n366) );
  NBUFFX2 U582 ( .IN(reset_n), .Q(n365) );
  NBUFFX2 U583 ( .IN(reset_n), .Q(n364) );
  NBUFFX2 U584 ( .IN(reset_n), .Q(n363) );
  NBUFFX2 U585 ( .IN(reset_n), .Q(n362) );
  NBUFFX2 U586 ( .IN(reset_n), .Q(n361) );
  XOR3X1 U587 ( .IN1(reg_b[13]), .IN2(reg_a[13]), .IN3(n467), .Q(n469) );
  OAI21X1 U588 ( .IN1(reg_a[13]), .IN2(n383), .IN3(n464), .QN(n471) );
  AO22X1 U589 ( .IN1(reg_a[13]), .IN2(n331), .IN3(result[13]), .IN4(n322), .Q(
        n73) );
  AO222X1 U590 ( .IN1(n268), .IN2(n155), .IN3(b_in[7]), .IN4(n149), .IN5(n154), 
        .IN6(n275), .Q(N99) );
  AO22X1 U591 ( .IN1(n155), .IN2(n342), .IN3(result[7]), .IN4(n306), .Q(n96)
         );
  INVX8 U592 ( .IN(n141), .QN(n233) );
  INVX8 U593 ( .IN(n141), .QN(n234) );
  INVX8 U594 ( .IN(n141), .QN(n602) );
  AO22X1 U595 ( .IN1(n242), .IN2(n343), .IN3(result[1]), .IN4(n307), .Q(n98)
         );
  OA21X1 U596 ( .IN1(n190), .IN2(n442), .IN3(n441), .Q(n443) );
  OA21X1 U597 ( .IN1(n571), .IN2(n172), .IN3(n570), .Q(n572) );
  NOR2X0 U598 ( .IN1(n592), .IN2(n591), .QN(n593) );
  NOR2X0 U599 ( .IN1(n531), .IN2(n591), .QN(n532) );
  AO222X1 U600 ( .IN1(n250), .IN2(n153), .IN3(b_in[2]), .IN4(n149), .IN5(
        reg_b[2]), .IN6(n275), .Q(N94) );
  OR4X1 U601 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n61) );
  AO221X1 U602 ( .IN1(n289), .IN2(n508), .IN3(a_in[22]), .IN4(n281), .IN5(n507), .Q(N81) );
  NBUFFX2 U603 ( .IN(n266), .Q(n265) );
  NBUFFX2 U604 ( .IN(n298), .Q(n258) );
  AO222X1 U605 ( .IN1(n256), .IN2(reg_a[30]), .IN3(b_in[30]), .IN4(n148), 
        .IN5(reg_b[30]), .IN6(n275), .Q(N122) );
  NBUFFX2 U606 ( .IN(n299), .Q(n256) );
  AO222X1 U607 ( .IN1(n254), .IN2(reg_a[24]), .IN3(b_in[24]), .IN4(n147), 
        .IN5(reg_b[24]), .IN6(n276), .Q(N116) );
  NBUFFX2 U608 ( .IN(n300), .Q(n254) );
  AO222X1 U609 ( .IN1(n261), .IN2(reg_a[19]), .IN3(b_in[19]), .IN4(n148), 
        .IN5(reg_b[19]), .IN6(n275), .Q(N111) );
  NBUFFX2 U610 ( .IN(n296), .Q(n261) );
  AO222X1 U611 ( .IN1(n264), .IN2(reg_a[12]), .IN3(b_in[12]), .IN4(n149), 
        .IN5(reg_b[12]), .IN6(n275), .Q(N104) );
  NBUFFX2 U612 ( .IN(n294), .Q(n264) );
  OR4X1 U613 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(
        reg_b[1]), .Q(n64) );
  NAND2X0 U614 ( .IN1(n527), .IN2(n526), .QN(n528) );
  AO22X1 U615 ( .IN1(n232), .IN2(n341), .IN3(result[5]), .IN4(n317), .Q(n94)
         );
  AO222X1 U616 ( .IN1(n263), .IN2(n237), .IN3(b_in[6]), .IN4(n147), .IN5(n113), 
        .IN6(n275), .Q(N98) );
  AO22X1 U617 ( .IN1(n237), .IN2(n342), .IN3(result[6]), .IN4(n317), .Q(n95)
         );
  AO222X1 U618 ( .IN1(n251), .IN2(n241), .IN3(b_in[4]), .IN4(n148), .IN5(n109), 
        .IN6(n275), .Q(N96) );
  XOR3X1 U619 ( .IN1(n241), .IN2(n109), .IN3(n571), .Q(n569) );
  AO22X1 U620 ( .IN1(n241), .IN2(n341), .IN3(result[4]), .IN4(n317), .Q(n93)
         );
  INVX2 U621 ( .IN(n244), .QN(n245) );
  AO221X1 U622 ( .IN1(n291), .IN2(n487), .IN3(a_in[17]), .IN4(n283), .IN5(n486), .Q(N76) );
  AO222X1 U623 ( .IN1(n266), .IN2(reg_a[9]), .IN3(b_in[9]), .IN4(n149), .IN5(
        reg_b[9]), .IN6(n276), .Q(N101) );
  AO222X1 U624 ( .IN1(n251), .IN2(reg_a[21]), .IN3(b_in[21]), .IN4(n147), 
        .IN5(reg_b[21]), .IN6(n275), .Q(N113) );
  AO222X1 U625 ( .IN1(n268), .IN2(reg_a[18]), .IN3(b_in[18]), .IN4(n149), 
        .IN5(reg_b[18]), .IN6(n276), .Q(N110) );
  AO222X1 U626 ( .IN1(n258), .IN2(reg_a[28]), .IN3(b_in[28]), .IN4(n149), 
        .IN5(reg_b[28]), .IN6(n275), .Q(N120) );
  AO222X1 U627 ( .IN1(n251), .IN2(n232), .IN3(b_in[5]), .IN4(n147), .IN5(n119), 
        .IN6(n276), .Q(N97) );
  AO222X1 U628 ( .IN1(n267), .IN2(n242), .IN3(b_in[1]), .IN4(n147), .IN5(
        reg_b[1]), .IN6(n276), .Q(N93) );
  AO222X1 U629 ( .IN1(n295), .IN2(reg_a[26]), .IN3(b_in[26]), .IN4(n147), 
        .IN5(reg_b[26]), .IN6(n275), .Q(N118) );
  AO222X1 U630 ( .IN1(n267), .IN2(reg_a[13]), .IN3(b_in[13]), .IN4(n147), 
        .IN5(reg_b[13]), .IN6(n276), .Q(N105) );
  AO222X1 U631 ( .IN1(n265), .IN2(n151), .IN3(b_in[8]), .IN4(n147), .IN5(n106), 
        .IN6(n276), .Q(N100) );
  NOR2X0 U632 ( .IN1(n159), .IN2(n239), .QN(n596) );
  AO221X1 U633 ( .IN1(n292), .IN2(n469), .IN3(a_in[13]), .IN4(n284), .IN5(n468), .Q(N72) );
  NBUFFX2 U634 ( .IN(n608), .Q(n250) );
  NBUFFX2 U635 ( .IN(n608), .Q(n251) );
  NBUFFX2 U636 ( .IN(n301), .Q(n252) );
  NBUFFX2 U637 ( .IN(n300), .Q(n253) );
  NBUFFX2 U638 ( .IN(n299), .Q(n255) );
  NBUFFX2 U639 ( .IN(n298), .Q(n257) );
  NBUFFX2 U640 ( .IN(n297), .Q(n259) );
  NBUFFX2 U641 ( .IN(n296), .Q(n260) );
  NBUFFX2 U642 ( .IN(n295), .Q(n262) );
  NBUFFX2 U643 ( .IN(n294), .Q(n263) );
  NBUFFX2 U644 ( .IN(n608), .Q(n300) );
  NBUFFX2 U645 ( .IN(n608), .Q(n299) );
  NBUFFX2 U646 ( .IN(n608), .Q(n298) );
  NBUFFX2 U647 ( .IN(n608), .Q(n297) );
  NBUFFX2 U648 ( .IN(n608), .Q(n296) );
  NBUFFX2 U649 ( .IN(n608), .Q(n295) );
  NBUFFX2 U650 ( .IN(n608), .Q(n294) );
  AND3X1 U651 ( .IN1(n376), .IN2(n272), .IN3(n134), .Q(n270) );
  NOR3X0 U652 ( .IN1(n270), .IN2(n501), .IN3(n413), .QN(n271) );
  NOR3X0 U653 ( .IN1(n412), .IN2(n497), .IN3(n498), .QN(n274) );
  AO221X1 U654 ( .IN1(n291), .IN2(n482), .IN3(a_in[16]), .IN4(n283), .IN5(n481), .Q(N75) );
  AO221X1 U655 ( .IN1(n288), .IN2(n544), .IN3(a_in[28]), .IN4(n280), .IN5(n543), .Q(N87) );
  AO221X1 U656 ( .IN1(n287), .IN2(n567), .IN3(a_in[3]), .IN4(n279), .IN5(n566), 
        .Q(N62) );
  AO22X1 U657 ( .IN1(n167), .IN2(reg_b[12]), .IN3(n233), .IN4(reg_a[12]), .Q(
        n462) );
  AO221X1 U658 ( .IN1(n290), .IN2(n500), .IN3(a_in[20]), .IN4(n282), .IN5(n499), .Q(N79) );
  AO22X1 U659 ( .IN1(n158), .IN2(reg_b[20]), .IN3(n602), .IN4(reg_a[20]), .Q(
        n499) );
  AO221X1 U660 ( .IN1(n291), .IN2(n474), .IN3(a_in[14]), .IN4(n283), .IN5(n473), .Q(N73) );
  AO22X1 U661 ( .IN1(n158), .IN2(reg_b[14]), .IN3(n234), .IN4(reg_a[14]), .Q(
        n473) );
  AO221X1 U662 ( .IN1(n292), .IN2(n460), .IN3(a_in[11]), .IN4(n284), .IN5(n459), .Q(N70) );
  AO22X1 U663 ( .IN1(n167), .IN2(reg_b[11]), .IN3(n602), .IN4(reg_a[11]), .Q(
        n459) );
  AO221X1 U664 ( .IN1(n290), .IN2(n495), .IN3(a_in[19]), .IN4(n282), .IN5(n494), .Q(N78) );
  AO22X1 U665 ( .IN1(n168), .IN2(reg_b[19]), .IN3(n602), .IN4(reg_a[19]), .Q(
        n494) );
  AO221X1 U666 ( .IN1(n290), .IN2(n503), .IN3(a_in[21]), .IN4(n282), .IN5(n502), .Q(N80) );
  AO22X1 U667 ( .IN1(n168), .IN2(reg_b[21]), .IN3(n234), .IN4(reg_a[21]), .Q(
        n502) );
  AO221X1 U668 ( .IN1(n290), .IN2(n490), .IN3(a_in[18]), .IN4(n282), .IN5(n489), .Q(N77) );
  AO22X1 U669 ( .IN1(n158), .IN2(reg_b[18]), .IN3(n602), .IN4(reg_a[18]), .Q(
        n489) );
  AO221X1 U670 ( .IN1(n291), .IN2(n477), .IN3(a_in[15]), .IN4(n283), .IN5(n476), .Q(N74) );
  AO22X1 U671 ( .IN1(n158), .IN2(reg_b[15]), .IN3(n233), .IN4(reg_a[15]), .Q(
        n476) );
  AO22X1 U672 ( .IN1(n167), .IN2(reg_b[0]), .IN3(n234), .IN4(reg_a[0]), .Q(
        n603) );
  AO22X1 U673 ( .IN1(n167), .IN2(reg_b[13]), .IN3(n234), .IN4(reg_a[13]), .Q(
        n468) );
  AO221X1 U674 ( .IN1(n292), .IN2(n454), .IN3(a_in[10]), .IN4(n284), .IN5(n453), .Q(N69) );
  AO22X1 U675 ( .IN1(n167), .IN2(reg_b[10]), .IN3(n233), .IN4(reg_a[10]), .Q(
        n453) );
  AO22X1 U676 ( .IN1(n167), .IN2(n109), .IN3(n602), .IN4(n241), .Q(n568) );
  OA21X1 U677 ( .IN1(n170), .IN2(n484), .IN3(n483), .Q(n485) );
  AO221X1 U678 ( .IN1(n287), .IN2(n569), .IN3(a_in[4]), .IN4(n279), .IN5(n568), 
        .Q(N63) );
  AO22X1 U679 ( .IN1(n168), .IN2(reg_b[31]), .IN3(n602), .IN4(reg_a[31]), .Q(
        n587) );
  AO221X1 U680 ( .IN1(n293), .IN2(n446), .IN3(a_in[8]), .IN4(n285), .IN5(n445), 
        .Q(N67) );
  AO22X1 U681 ( .IN1(n168), .IN2(n106), .IN3(n233), .IN4(n151), .Q(n445) );
  AO221X1 U682 ( .IN1(n288), .IN2(n541), .IN3(a_in[27]), .IN4(n280), .IN5(n540), .Q(N86) );
  AO22X1 U683 ( .IN1(n158), .IN2(reg_b[27]), .IN3(n233), .IN4(reg_a[27]), .Q(
        n540) );
  AO221X1 U684 ( .IN1(n288), .IN2(n551), .IN3(a_in[29]), .IN4(n280), .IN5(n550), .Q(N88) );
  AO22X1 U685 ( .IN1(n167), .IN2(reg_b[29]), .IN3(n234), .IN4(reg_a[29]), .Q(
        n550) );
  AO221X1 U686 ( .IN1(n286), .IN2(n583), .IN3(a_in[7]), .IN4(n278), .IN5(n582), 
        .Q(N66) );
  AO22X1 U687 ( .IN1(n168), .IN2(n154), .IN3(n602), .IN4(n155), .Q(n582) );
  AO221X1 U688 ( .IN1(n287), .IN2(n561), .IN3(a_in[2]), .IN4(n279), .IN5(n560), 
        .Q(N61) );
  AO22X1 U689 ( .IN1(n167), .IN2(reg_b[2]), .IN3(n602), .IN4(n153), .Q(n560)
         );
  AO221X1 U690 ( .IN1(n289), .IN2(n523), .IN3(a_in[25]), .IN4(n281), .IN5(n522), .Q(N84) );
  AO22X1 U691 ( .IN1(n168), .IN2(reg_b[25]), .IN3(n233), .IN4(reg_a[25]), .Q(
        n522) );
  AO22X1 U692 ( .IN1(n158), .IN2(reg_b[16]), .IN3(n602), .IN4(reg_a[16]), .Q(
        n481) );
  AO22X1 U693 ( .IN1(n158), .IN2(reg_b[17]), .IN3(n233), .IN4(n103), .Q(n486)
         );
  AO22X1 U694 ( .IN1(n168), .IN2(n119), .IN3(n234), .IN4(n232), .Q(n573) );
  OA21X1 U695 ( .IN1(n171), .IN2(n471), .IN3(n470), .Q(n472) );
  AO221X1 U696 ( .IN1(n289), .IN2(n513), .IN3(a_in[23]), .IN4(n281), .IN5(n512), .Q(N82) );
  AO22X1 U697 ( .IN1(n158), .IN2(reg_b[23]), .IN3(n234), .IN4(reg_a[23]), .Q(
        n512) );
  AO221X1 U698 ( .IN1(n287), .IN2(n574), .IN3(a_in[5]), .IN4(n279), .IN5(n573), 
        .Q(N64) );
  AO222X1 U699 ( .IN1(reg_a[0]), .IN2(n267), .IN3(b_in[0]), .IN4(n149), .IN5(
        reg_b[0]), .IN6(n276), .Q(N92) );
  OR4X1 U700 ( .IN1(reg_b[0]), .IN2(reg_b[10]), .IN3(reg_b[11]), .IN4(
        reg_b[12]), .Q(n66) );
  AO221X1 U701 ( .IN1(n286), .IN2(n577), .IN3(a_in[6]), .IN4(n278), .IN5(n576), 
        .Q(N65) );
  AO22X1 U702 ( .IN1(n168), .IN2(n113), .IN3(n233), .IN4(n237), .Q(n576) );
  AO221X1 U703 ( .IN1(n289), .IN2(n517), .IN3(a_in[24]), .IN4(n281), .IN5(n516), .Q(N83) );
  AO22X1 U704 ( .IN1(n158), .IN2(reg_b[24]), .IN3(n234), .IN4(reg_a[24]), .Q(
        n516) );
  AO22X1 U705 ( .IN1(n158), .IN2(reg_b[22]), .IN3(n602), .IN4(reg_a[22]), .Q(
        n507) );
  AO221X1 U706 ( .IN1(n293), .IN2(n449), .IN3(a_in[9]), .IN4(n285), .IN5(n448), 
        .Q(N68) );
  AO22X1 U707 ( .IN1(n167), .IN2(reg_b[9]), .IN3(n234), .IN4(reg_a[9]), .Q(
        n448) );
  AO221X1 U708 ( .IN1(n292), .IN2(n463), .IN3(a_in[12]), .IN4(n284), .IN5(n462), .Q(N71) );
  OA21X1 U709 ( .IN1(n124), .IN2(n456), .IN3(n455), .Q(n458) );
  AO221X1 U710 ( .IN1(n286), .IN2(n605), .IN3(a_in[0]), .IN4(n278), .IN5(n603), 
        .Q(N59) );
  AO221X1 U711 ( .IN1(n588), .IN2(n286), .IN3(a_in[31]), .IN4(n278), .IN5(n587), .Q(N90) );
  AO22X1 U712 ( .IN1(n158), .IN2(reg_b[28]), .IN3(n233), .IN4(reg_a[28]), .Q(
        n543) );
  NBUFFX2 U713 ( .IN(n608), .Q(n301) );
  AO22X1 U714 ( .IN1(n168), .IN2(reg_b[3]), .IN3(n233), .IN4(reg_a[3]), .Q(
        n566) );
  INVX4 U715 ( .IN(n539), .QN(n420) );
  OR2X2 U716 ( .IN1(n245), .IN2(n273), .Q(n601) );
  NOR2X4 U717 ( .IN1(n419), .IN2(n418), .QN(n539) );
  NAND2X4 U718 ( .IN1(n420), .IN2(n421), .QN(n422) );
  NAND2X4 U719 ( .IN1(n165), .IN2(n424), .QN(n425) );
  NAND2X4 U720 ( .IN1(n426), .IN2(n425), .QN(n547) );
  NOR2X4 U721 ( .IN1(n547), .IN2(n427), .QN(n428) );
  NAND2X4 U722 ( .IN1(n429), .IN2(n430), .QN(n431) );
  INVX8 U723 ( .IN(n590), .QN(n604) );
endmodule

