module fifo (	
	 input            wr_clk,   //write clock
         input            rd_clk,   //read clock
         input            reset_n,  //reset async active low
         input            wr,       //write enable 
         input            rd,       //read enable    
         input      [7:0] data_in,  //data in
         output reg [7:0] data_out, //data out
         output           empty,    //empty flag
         output           full      //full flag
        );

    


endmodule
