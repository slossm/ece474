
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, n6, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ns;

  DFFARX1 \reg_b_reg[0]  ( .D(N92), .CLK(clk), .RSTB(n377), .Q(reg_b[0]), .QN(
        n307) );
  DFFARX1 \reg_b_reg[1]  ( .D(N93), .CLK(clk), .RSTB(n377), .Q(reg_b[1]), .QN(
        n297) );
  DFFARX1 \reg_b_reg[4]  ( .D(N96), .CLK(clk), .RSTB(n374), .QN(n134) );
  DFFARX1 \gcd_ps_reg[0]  ( .D(gcd_ns[0]), .CLK(clk), .RSTB(n378), .Q(n264), 
        .QN(n67) );
  DFFARX1 \reg_a_reg[20]  ( .D(N79), .CLK(clk), .RSTB(n368), .Q(reg_a[20]), 
        .QN(n236) );
  DFFARX1 \reg_a_reg[11]  ( .D(N70), .CLK(clk), .RSTB(n363), .Q(reg_a[11]), 
        .QN(n194) );
  DFFARX1 \gcd_ps_reg[1]  ( .D(gcd_ns[1]), .CLK(clk), .RSTB(n377), .Q(n282), 
        .QN(n100) );
  DFFARX1 \reg_b_reg[29]  ( .D(N121), .CLK(clk), .RSTB(n372), .Q(reg_b[29]), 
        .QN(n274) );
  DFFARX1 \reg_b_reg[30]  ( .D(N122), .CLK(clk), .RSTB(n373), .Q(reg_b[30]), 
        .QN(n275) );
  DFFARX1 \reg_b_reg[11]  ( .D(N103), .CLK(clk), .RSTB(n363), .Q(reg_b[11]), 
        .QN(n191) );
  DFFARX1 \reg_a_reg[19]  ( .D(N78), .CLK(clk), .RSTB(n367), .Q(reg_a[19]), 
        .QN(n234) );
  DFFARX1 \reg_a_reg[16]  ( .D(N75), .CLK(clk), .RSTB(n366), .Q(reg_a[16]), 
        .QN(n241) );
  DFFARX1 \reg_a_reg[18]  ( .D(N77), .CLK(clk), .RSTB(n367), .Q(reg_a[18]), 
        .QN(n271) );
  DFFARX1 \reg_b_reg[25]  ( .D(N117), .CLK(clk), .RSTB(n370), .Q(reg_b[25]), 
        .QN(n278) );
  DFFARX1 \reg_b_reg[21]  ( .D(N113), .CLK(clk), .RSTB(n368), .Q(reg_b[21]), 
        .QN(n279) );
  DFFARX1 \reg_b_reg[10]  ( .D(N102), .CLK(clk), .RSTB(n363), .Q(reg_b[10]), 
        .QN(n277) );
  DFFARX1 \reg_b_reg[18]  ( .D(N110), .CLK(clk), .RSTB(n367), .Q(reg_b[18]), 
        .QN(n266) );
  DFFARX1 \reg_b_reg[22]  ( .D(N114), .CLK(clk), .RSTB(n369), .Q(reg_b[22]), 
        .QN(n281) );
  DFFARX1 \reg_b_reg[24]  ( .D(N116), .CLK(clk), .RSTB(n370), .Q(reg_b[24]), 
        .QN(n269) );
  DFFARX1 \reg_b_reg[19]  ( .D(N111), .CLK(clk), .RSTB(n367), .Q(reg_b[19]), 
        .QN(n268) );
  DFFARX1 \reg_b_reg[15]  ( .D(N107), .CLK(clk), .RSTB(n365), .Q(reg_b[15]), 
        .QN(n265) );
  DFFARX1 \reg_b_reg[16]  ( .D(N108), .CLK(clk), .RSTB(n366), .Q(reg_b[16]), 
        .QN(n232) );
  DFFARX1 \reg_b_reg[9]  ( .D(N101), .CLK(clk), .RSTB(n362), .Q(reg_b[9]), 
        .QN(n280) );
  DFFARX1 \reg_b_reg[12]  ( .D(N104), .CLK(clk), .RSTB(n364), .Q(reg_b[12]), 
        .QN(n267) );
  DFFARX1 \reg_a_reg[31]  ( .D(N90), .CLK(clk), .RSTB(n376), .Q(reg_a[31]), 
        .QN(n230) );
  DFFARX1 \reg_b_reg[2]  ( .D(N94), .CLK(clk), .RSTB(n373), .Q(reg_b[2]), .QN(
        n262) );
  DFFARX1 \reg_b_reg[8]  ( .D(N100), .CLK(clk), .RSTB(n362), .Q(reg_b[8]), 
        .QN(n202) );
  DFFARX1 \reg_a_reg[2]  ( .D(N61), .CLK(clk), .RSTB(n373), .Q(reg_a[2]), .QN(
        n260) );
  DFFARX1 \reg_a_reg[7]  ( .D(N66), .CLK(clk), .RSTB(n376), .QN(n199) );
  DFFARX1 \reg_a_reg[4]  ( .D(N63), .CLK(clk), .RSTB(n374), .QN(n289) );
  DFFARX1 \reg_a_reg[9]  ( .D(N68), .CLK(clk), .RSTB(n362), .Q(reg_a[9]), .QN(
        n135) );
  DFFARX1 \reg_a_reg[6]  ( .D(N65), .CLK(clk), .RSTB(n375), .Q(n196), .QN(n215) );
  DFFARX1 \result_reg[31]  ( .D(n97), .CLK(clk), .RSTB(n376), .Q(result[31])
         );
  DFFARX1 \result_reg[7]  ( .D(n96), .CLK(clk), .RSTB(n376), .Q(result[7]) );
  DFFARX1 \result_reg[1]  ( .D(n98), .CLK(clk), .RSTB(n377), .Q(result[1]) );
  DFFARX1 \result_reg[8]  ( .D(n68), .CLK(clk), .RSTB(n362), .Q(result[8]) );
  DFFARX1 \result_reg[20]  ( .D(n80), .CLK(clk), .RSTB(n368), .Q(result[20])
         );
  DFFARX1 \result_reg[19]  ( .D(n79), .CLK(clk), .RSTB(n367), .Q(result[19])
         );
  DFFARX1 \result_reg[18]  ( .D(n78), .CLK(clk), .RSTB(n367), .Q(result[18])
         );
  DFFARX1 \result_reg[17]  ( .D(n77), .CLK(clk), .RSTB(n366), .Q(result[17])
         );
  DFFARX1 \result_reg[16]  ( .D(n76), .CLK(clk), .RSTB(n366), .Q(result[16])
         );
  DFFARX1 \result_reg[15]  ( .D(n75), .CLK(clk), .RSTB(n365), .Q(result[15])
         );
  DFFARX1 \result_reg[14]  ( .D(n74), .CLK(clk), .RSTB(n365), .Q(result[14])
         );
  DFFARX1 \result_reg[13]  ( .D(n73), .CLK(clk), .RSTB(n364), .Q(result[13])
         );
  DFFARX1 \result_reg[12]  ( .D(n72), .CLK(clk), .RSTB(n364), .Q(result[12])
         );
  DFFARX1 \result_reg[11]  ( .D(n71), .CLK(clk), .RSTB(n363), .Q(result[11])
         );
  DFFARX1 \result_reg[10]  ( .D(n70), .CLK(clk), .RSTB(n363), .Q(result[10])
         );
  DFFARX1 \result_reg[9]  ( .D(n69), .CLK(clk), .RSTB(n362), .Q(result[9]) );
  DFFARX1 \result_reg[30]  ( .D(n90), .CLK(clk), .RSTB(n373), .Q(result[30])
         );
  DFFARX1 \result_reg[29]  ( .D(n89), .CLK(clk), .RSTB(n372), .Q(result[29])
         );
  DFFARX1 \result_reg[28]  ( .D(n88), .CLK(clk), .RSTB(n372), .Q(result[28])
         );
  DFFARX1 \result_reg[27]  ( .D(n87), .CLK(clk), .RSTB(n371), .Q(result[27])
         );
  DFFARX1 \result_reg[26]  ( .D(n86), .CLK(clk), .RSTB(n371), .Q(result[26])
         );
  DFFARX1 \result_reg[25]  ( .D(n85), .CLK(clk), .RSTB(n370), .Q(result[25])
         );
  DFFARX1 \result_reg[24]  ( .D(n84), .CLK(clk), .RSTB(n370), .Q(result[24])
         );
  DFFARX1 \result_reg[23]  ( .D(n83), .CLK(clk), .RSTB(n369), .Q(result[23])
         );
  DFFARX1 \result_reg[22]  ( .D(n82), .CLK(clk), .RSTB(n369), .Q(result[22])
         );
  DFFARX1 \result_reg[21]  ( .D(n81), .CLK(clk), .RSTB(n368), .Q(result[21])
         );
  DFFARX1 \result_reg[6]  ( .D(n95), .CLK(clk), .RSTB(n375), .Q(result[6]) );
  DFFARX1 \result_reg[5]  ( .D(n94), .CLK(clk), .RSTB(n375), .Q(result[5]) );
  DFFARX1 \result_reg[4]  ( .D(n93), .CLK(clk), .RSTB(n374), .Q(result[4]) );
  DFFARX1 \result_reg[3]  ( .D(n92), .CLK(clk), .RSTB(n374), .Q(result[3]) );
  DFFARX1 \result_reg[2]  ( .D(n91), .CLK(clk), .RSTB(n373), .Q(result[2]) );
  DFFARX1 \result_reg[0]  ( .D(n99), .CLK(clk), .RSTB(n377), .Q(result[0]) );
  DFFARX1 \reg_a_reg[26]  ( .D(N85), .CLK(clk), .RSTB(n371), .Q(reg_a[26]), 
        .QN(n546) );
  DFFARX1 \reg_b_reg[3]  ( .D(N95), .CLK(clk), .RSTB(n374), .Q(reg_b[3]) );
  DFFARX1 \reg_b_reg[27]  ( .D(N119), .CLK(clk), .RSTB(n371), .Q(reg_b[27]) );
  DFFARX1 \reg_b_reg[14]  ( .D(N106), .CLK(clk), .RSTB(n365), .Q(reg_b[14]), 
        .QN(n398) );
  DFFARX1 \reg_b_reg[31]  ( .D(N123), .CLK(clk), .RSTB(n376), .Q(reg_b[31]), 
        .QN(n595) );
  DFFARX1 \reg_b_reg[20]  ( .D(N112), .CLK(clk), .RSTB(n368), .Q(reg_b[20]), 
        .QN(n392) );
  DFFARX1 \reg_b_reg[28]  ( .D(N120), .CLK(clk), .RSTB(n372), .Q(reg_b[28]) );
  DFFARX1 \reg_b_reg[13]  ( .D(N105), .CLK(clk), .RSTB(n364), .Q(reg_b[13]), 
        .QN(n401) );
  DFFARX1 \reg_b_reg[23]  ( .D(N115), .CLK(clk), .RSTB(n369), .Q(reg_b[23]), 
        .QN(n389) );
  DFFARX1 \reg_b_reg[17]  ( .D(N109), .CLK(clk), .RSTB(n366), .Q(reg_b[17]), 
        .QN(n395) );
  DFFARX1 \reg_b_reg[26]  ( .D(N118), .CLK(clk), .RSTB(n371), .Q(reg_b[26]), 
        .QN(n388) );
  DFFARX1 \reg_a_reg[30]  ( .D(N89), .CLK(clk), .RSTB(n373), .Q(reg_a[30]) );
  DFFARX1 \reg_a_reg[29]  ( .D(N88), .CLK(clk), .RSTB(n372), .Q(reg_a[29]) );
  DFFARX1 \reg_a_reg[25]  ( .D(N84), .CLK(clk), .RSTB(n370), .Q(reg_a[25]) );
  DFFARX1 \reg_a_reg[14]  ( .D(N73), .CLK(clk), .RSTB(n365), .Q(reg_a[14]) );
  DFFARX1 \reg_a_reg[23]  ( .D(N82), .CLK(clk), .RSTB(n369), .Q(reg_a[23]) );
  DFFARX1 \reg_a_reg[17]  ( .D(N76), .CLK(clk), .RSTB(n366), .Q(reg_a[17]) );
  DFFARX1 \reg_a_reg[27]  ( .D(N86), .CLK(clk), .RSTB(n371), .Q(reg_a[27]), 
        .QN(n442) );
  DFFARX1 \reg_a_reg[22]  ( .D(N81), .CLK(clk), .RSTB(n369), .Q(reg_a[22]) );
  DFFARX1 \reg_b_reg[5]  ( .D(N97), .CLK(clk), .RSTB(n375), .QN(n292) );
  DFFARX1 \reg_b_reg[6]  ( .D(N98), .CLK(clk), .RSTB(n375), .QN(n287) );
  DFFARX1 \reg_b_reg[7]  ( .D(N99), .CLK(clk), .RSTB(n376), .QN(n261) );
  DFFARX1 \reg_a_reg[13]  ( .D(N72), .CLK(clk), .RSTB(n364), .Q(reg_a[13]), 
        .QN(n240) );
  DFFARX1 \reg_a_reg[3]  ( .D(N62), .CLK(clk), .RSTB(n374), .Q(reg_a[3]), .QN(
        n239) );
  DFFARX1 \reg_a_reg[28]  ( .D(N87), .CLK(clk), .RSTB(n372), .Q(reg_a[28]), 
        .QN(n263) );
  DFFARX1 \reg_a_reg[15]  ( .D(N74), .CLK(clk), .RSTB(n365), .Q(reg_a[15]), 
        .QN(n272) );
  DFFARX1 \reg_a_reg[24]  ( .D(N83), .CLK(clk), .RSTB(n370), .Q(reg_a[24]), 
        .QN(n270) );
  DFFARX1 \reg_a_reg[12]  ( .D(N71), .CLK(clk), .RSTB(n364), .Q(reg_a[12]), 
        .QN(n276) );
  DFFARX1 \reg_a_reg[21]  ( .D(N80), .CLK(clk), .RSTB(n368), .Q(reg_a[21]), 
        .QN(n273) );
  DFFARX1 \reg_a_reg[0]  ( .D(N59), .CLK(clk), .RSTB(n378), .Q(reg_a[0]), .QN(
        n298) );
  DFFARX1 \reg_a_reg[5]  ( .D(N64), .CLK(clk), .RSTB(n375), .QN(n197) );
  DFFARX1 \reg_a_reg[10]  ( .D(N69), .CLK(clk), .RSTB(n363), .Q(reg_a[10]), 
        .QN(n192) );
  DFFARX1 \reg_a_reg[8]  ( .D(N67), .CLK(clk), .RSTB(n362), .Q(reg_a[8]), .QN(
        n200) );
  DFFARX2 \reg_a_reg[1]  ( .D(N60), .CLK(clk), .RSTB(n377), .QN(n211) );
  NAND2X4 U166 ( .IN1(n189), .IN2(n443), .QN(n444) );
  NAND2X4 U167 ( .IN1(n441), .IN2(n190), .QN(n189) );
  NBUFFX16 U168 ( .IN(reg_b[3]), .Q(n102) );
  NAND2X4 U169 ( .IN1(n212), .IN2(n608), .QN(n213) );
  NAND2X4 U170 ( .IN1(n448), .IN2(n449), .QN(n450) );
  NOR2X4 U171 ( .IN1(n408), .IN2(n407), .QN(n409) );
  NOR2X1 U172 ( .IN1(n406), .IN2(n405), .QN(n408) );
  INVX4 U173 ( .IN(n205), .QN(n103) );
  INVX4 U174 ( .IN(n205), .QN(n104) );
  INVX2 U175 ( .IN(n302), .QN(n303) );
  INVX4 U176 ( .IN(n205), .QN(n615) );
  OR2X2 U177 ( .IN1(n608), .IN2(n455), .Q(n302) );
  OR2X2 U178 ( .IN1(n608), .IN2(n455), .Q(n205) );
  NAND2X1 U179 ( .IN1(n262), .IN2(n198), .QN(n573) );
  NOR2X1 U180 ( .IN1(n211), .IN2(n291), .QN(n605) );
  NAND2X2 U181 ( .IN1(n211), .IN2(n209), .QN(n210) );
  INVX4 U182 ( .IN(n211), .QN(n296) );
  NAND2X4 U183 ( .IN1(n470), .IN2(n421), .QN(n422) );
  INVX2 U184 ( .IN(n466), .QN(n421) );
  NOR2X4 U185 ( .IN1(n412), .IN2(n461), .QN(n214) );
  INVX1 U186 ( .IN(n414), .QN(n404) );
  OR2X2 U187 ( .IN1(n284), .IN2(n292), .Q(n414) );
  NBUFFX2 U188 ( .IN(n310), .Q(n105) );
  NBUFFX8 U189 ( .IN(n310), .Q(n106) );
  NBUFFX16 U190 ( .IN(n310), .Q(n107) );
  INVX2 U191 ( .IN(n312), .QN(n310) );
  INVX0 U192 ( .IN(n528), .QN(n187) );
  OR2X1 U193 ( .IN1(reg_a[17]), .IN2(n395), .Q(n397) );
  INVX0 U194 ( .IN(n524), .QN(n390) );
  OR2X1 U195 ( .IN1(reg_a[14]), .IN2(n398), .Q(n400) );
  NAND2X2 U196 ( .IN1(n415), .IN2(n414), .QN(n207) );
  OR2X2 U197 ( .IN1(n404), .IN2(n228), .Q(n458) );
  INVX0 U198 ( .IN(n403), .QN(n424) );
  NAND2X0 U199 ( .IN1(n276), .IN2(reg_b[12]), .QN(n483) );
  INVX0 U200 ( .IN(n397), .QN(n428) );
  INVX0 U201 ( .IN(n500), .QN(n396) );
  NOR4X0 U202 ( .IN1(n61), .IN2(n62), .IN3(n59), .IN4(n60), .QN(n243) );
  NOR4X0 U203 ( .IN1(n65), .IN2(n66), .IN3(n63), .IN4(n64), .QN(n242) );
  INVX4 U204 ( .IN(n216), .QN(n286) );
  INVX4 U205 ( .IN(n217), .QN(n285) );
  NAND2X0 U206 ( .IN1(n277), .IN2(n193), .QN(n474) );
  INVX0 U207 ( .IN(n192), .QN(n193) );
  NAND2X2 U208 ( .IN1(n430), .IN2(n133), .QN(n301) );
  INVX0 U209 ( .IN(n514), .QN(n306) );
  NOR2X0 U210 ( .IN1(n404), .IN2(n228), .QN(n218) );
  OR2X1 U211 ( .IN1(reg_a[20]), .IN2(n392), .Q(n394) );
  NOR2X0 U212 ( .IN1(n537), .IN2(n111), .QN(n434) );
  AO22X1 U213 ( .IN1(n393), .IN2(n394), .IN3(reg_a[20]), .IN4(n392), .Q(n517)
         );
  INVX0 U214 ( .IN(n513), .QN(n393) );
  NAND2X0 U215 ( .IN1(n270), .IN2(reg_b[24]), .QN(n531) );
  OR4X1 U216 ( .IN1(reg_b[0]), .IN2(reg_b[10]), .IN3(reg_b[11]), .IN4(
        reg_b[12]), .Q(n66) );
  INVX0 U217 ( .IN(n419), .QN(n412) );
  INVX0 U218 ( .IN(n433), .QN(n529) );
  NAND2X0 U219 ( .IN1(n267), .IN2(reg_a[12]), .QN(n484) );
  NAND2X2 U220 ( .IN1(n210), .IN2(n610), .QN(n568) );
  INVX0 U221 ( .IN(n297), .QN(n209) );
  NAND2X1 U222 ( .IN1(n297), .IN2(n296), .QN(n569) );
  AND2X1 U223 ( .IN1(n445), .IN2(n444), .Q(n148) );
  NAND2X0 U224 ( .IN1(n272), .IN2(reg_b[15]), .QN(n495) );
  NAND2X0 U225 ( .IN1(n271), .IN2(reg_b[18]), .QN(n508) );
  OAI21X1 U226 ( .IN1(reg_a[19]), .IN2(n268), .IN3(n508), .QN(n514) );
  NAND2X0 U227 ( .IN1(n268), .IN2(reg_a[19]), .QN(n513) );
  INVX0 U228 ( .IN(n430), .QN(n515) );
  NBUFFX2 U229 ( .IN(n226), .Q(n139) );
  XOR3X1 U230 ( .IN1(reg_b[14]), .IN2(reg_a[14]), .IN3(n490), .Q(n491) );
  NBUFFX2 U231 ( .IN(n227), .Q(n183) );
  XOR3X1 U232 ( .IN1(reg_a[9]), .IN2(reg_b[9]), .IN3(n254), .Q(n468) );
  XOR3X1 U233 ( .IN1(reg_b[8]), .IN2(reg_a[8]), .IN3(n462), .Q(n465) );
  XOR3X1 U234 ( .IN1(n284), .IN2(n293), .IN3(n582), .Q(n583) );
  INVX2 U235 ( .IN(n197), .QN(n284) );
  NBUFFX2 U236 ( .IN(n251), .Q(n184) );
  AND2X1 U237 ( .IN1(n568), .IN2(n569), .Q(n253) );
  NBUFFX2 U238 ( .IN(n612), .Q(n314) );
  OA21X1 U239 ( .IN1(n148), .IN2(n564), .IN3(n563), .Q(n248) );
  NAND2X0 U240 ( .IN1(n265), .IN2(reg_a[15]), .QN(n496) );
  NBUFFX2 U241 ( .IN(n252), .Q(n222) );
  NBUFFX2 U242 ( .IN(n612), .Q(n317) );
  NAND2X0 U243 ( .IN1(n266), .IN2(reg_a[18]), .QN(n509) );
  NBUFFX2 U244 ( .IN(n225), .Q(n138) );
  INVX2 U245 ( .IN(n289), .QN(n294) );
  XOR3X1 U246 ( .IN1(reg_b[27]), .IN2(reg_a[27]), .IN3(n551), .Q(n553) );
  NAND2X1 U247 ( .IN1(n119), .IN2(n155), .QN(N82) );
  XOR3X1 U248 ( .IN1(n288), .IN2(n295), .IN3(n247), .Q(n586) );
  XOR3X1 U249 ( .IN1(n203), .IN2(n204), .IN3(n590), .Q(n592) );
  XOR3X1 U250 ( .IN1(reg_b[28]), .IN2(reg_a[28]), .IN3(n149), .Q(n555) );
  AND2X1 U251 ( .IN1(n441), .IN2(n190), .Q(n149) );
  NAND2X0 U252 ( .IN1(n607), .IN2(n606), .QN(N60) );
  NOR2X0 U253 ( .IN1(n605), .IN2(n604), .QN(n606) );
  INVX0 U254 ( .IN(n158), .QN(n159) );
  INVX0 U255 ( .IN(n608), .QN(n158) );
  XOR3X1 U256 ( .IN1(reg_b[11]), .IN2(reg_a[11]), .IN3(n477), .Q(n479) );
  NAND3X0 U257 ( .IN1(n433), .IN2(n187), .IN3(n532), .QN(n108) );
  NAND2X4 U258 ( .IN1(n450), .IN2(n451), .QN(n109) );
  NOR2X0 U259 ( .IN1(reg_a[30]), .IN2(n275), .QN(n110) );
  NOR2X0 U260 ( .IN1(reg_a[26]), .IN2(n388), .QN(n111) );
  AND2X1 U261 ( .IN1(n249), .IN2(n391), .Q(n112) );
  INVX0 U262 ( .IN(n292), .QN(n293) );
  AND2X1 U263 ( .IN1(n300), .IN2(n520), .Q(n113) );
  OR2X1 U264 ( .IN1(n489), .IN2(n426), .Q(n114) );
  NOR2X0 U265 ( .IN1(n456), .IN2(n259), .QN(n115) );
  OR2X1 U266 ( .IN1(n501), .IN2(n428), .Q(n116) );
  NAND2X0 U267 ( .IN1(n242), .IN2(n243), .QN(n6) );
  OR2X1 U268 ( .IN1(n480), .IN2(n425), .Q(n117) );
  OR2X1 U269 ( .IN1(n492), .IN2(n427), .Q(n118) );
  NBUFFX2 U270 ( .IN(n612), .Q(n316) );
  NBUFFX8 U271 ( .IN(n612), .Q(n313) );
  AOI22X1 U272 ( .IN1(n223), .IN2(reg_b[23]), .IN3(n286), .IN4(reg_a[23]), 
        .QN(n119) );
  OR2X1 U273 ( .IN1(n212), .IN2(n283), .Q(n454) );
  AOI22X1 U274 ( .IN1(n221), .IN2(reg_b[25]), .IN3(n285), .IN4(reg_a[25]), 
        .QN(n120) );
  AOI22X1 U275 ( .IN1(n223), .IN2(reg_b[29]), .IN3(n286), .IN4(reg_a[29]), 
        .QN(n121) );
  AOI22X1 U276 ( .IN1(n220), .IN2(reg_b[30]), .IN3(n286), .IN4(reg_a[30]), 
        .QN(n122) );
  AOI22X1 U277 ( .IN1(n224), .IN2(reg_b[9]), .IN3(n286), .IN4(reg_a[9]), .QN(
        n123) );
  AOI22X1 U278 ( .IN1(n220), .IN2(reg_b[14]), .IN3(n286), .IN4(reg_a[14]), 
        .QN(n124) );
  AOI22X1 U279 ( .IN1(n220), .IN2(reg_b[24]), .IN3(n286), .IN4(reg_a[24]), 
        .QN(n125) );
  AOI22X1 U280 ( .IN1(n220), .IN2(reg_b[13]), .IN3(n161), .IN4(reg_a[13]), 
        .QN(n126) );
  AOI22X1 U281 ( .IN1(n221), .IN2(reg_b[20]), .IN3(n161), .IN4(reg_a[20]), 
        .QN(n127) );
  AOI22X1 U282 ( .IN1(n221), .IN2(reg_b[21]), .IN3(n286), .IN4(reg_a[21]), 
        .QN(n128) );
  AOI22X1 U283 ( .IN1(n224), .IN2(reg_b[8]), .IN3(n286), .IN4(reg_a[8]), .QN(
        n129) );
  AOI22X1 U284 ( .IN1(n221), .IN2(n293), .IN3(n286), .IN4(n284), .QN(n130) );
  AOI22X1 U285 ( .IN1(n224), .IN2(reg_b[0]), .IN3(n286), .IN4(reg_a[0]), .QN(
        n131) );
  INVX2 U286 ( .IN(n261), .QN(n203) );
  OR2X1 U287 ( .IN1(n475), .IN2(n424), .Q(n132) );
  INVX2 U288 ( .IN(n134), .QN(n290) );
  AND2X1 U289 ( .IN1(n306), .IN2(n394), .Q(n133) );
  NAND2X0 U290 ( .IN1(n264), .IN2(n100), .QN(n455) );
  INVX0 U291 ( .IN(n196), .QN(n413) );
  NAND2X2 U292 ( .IN1(n214), .IN2(n459), .QN(n417) );
  OR2X1 U293 ( .IN1(n416), .IN2(n584), .Q(n459) );
  IBUFFX2 U294 ( .IN(n464), .QN(n245) );
  NAND2X4 U295 ( .IN1(n135), .IN2(reg_b[9]), .QN(n469) );
  NOR2X4 U296 ( .IN1(n455), .IN2(n452), .QN(n147) );
  INVX8 U297 ( .IN(n156), .QN(n136) );
  INVX8 U298 ( .IN(n156), .QN(n137) );
  NAND2X0 U299 ( .IN1(n103), .IN2(n288), .QN(n140) );
  NAND2X0 U300 ( .IN1(b_in[6]), .IN2(n137), .QN(n141) );
  NAND2X0 U301 ( .IN1(n295), .IN2(n107), .QN(n142) );
  NAND3X0 U302 ( .IN1(n140), .IN2(n141), .IN3(n142), .QN(N98) );
  OAI21X2 U303 ( .IN1(reg_a[10]), .IN2(n277), .IN3(n469), .QN(n475) );
  NAND2X2 U304 ( .IN1(n105), .IN2(n245), .QN(n291) );
  NAND2X2 U305 ( .IN1(n452), .IN2(n212), .QN(n453) );
  NAND2X0 U306 ( .IN1(n614), .IN2(n516), .QN(n143) );
  NAND2X0 U307 ( .IN1(a_in[20]), .IN2(n316), .QN(n144) );
  NAND3X0 U308 ( .IN1(n143), .IN2(n144), .IN3(n127), .QN(N79) );
  NAND2X2 U309 ( .IN1(n145), .IN2(n203), .QN(n146) );
  NAND2X2 U310 ( .IN1(n146), .IN2(n587), .QN(n461) );
  INVX0 U311 ( .IN(n204), .QN(n145) );
  NOR2X4 U312 ( .IN1(n147), .IN2(n456), .QN(n157) );
  INVX4 U313 ( .IN(n199), .QN(n204) );
  OR2X1 U314 ( .IN1(n288), .IN2(n287), .Q(n587) );
  OR2X1 U315 ( .IN1(n412), .IN2(n461), .Q(n467) );
  INVX8 U316 ( .IN(n157), .QN(n188) );
  INVX8 U317 ( .IN(n109), .QN(n608) );
  OR2X1 U318 ( .IN1(n263), .IN2(reg_b[28]), .Q(n445) );
  NAND2X0 U319 ( .IN1(n614), .IN2(n535), .QN(n150) );
  NAND2X0 U320 ( .IN1(a_in[25]), .IN2(n313), .QN(n151) );
  NAND3X0 U321 ( .IN1(n150), .IN2(n151), .IN3(n120), .QN(N84) );
  NAND2X0 U322 ( .IN1(n614), .IN2(n487), .QN(n152) );
  NAND2X0 U323 ( .IN1(a_in[13]), .IN2(n318), .QN(n153) );
  NAND3X0 U324 ( .IN1(n152), .IN2(n153), .IN3(n126), .QN(N72) );
  NBUFFX16 U325 ( .IN(n612), .Q(n318) );
  NOR2X4 U326 ( .IN1(n312), .IN2(n464), .QN(n206) );
  NAND2X1 U327 ( .IN1(n609), .IN2(n463), .QN(n216) );
  NAND2X2 U328 ( .IN1(n181), .IN2(n180), .QN(n154) );
  INVX2 U329 ( .IN(n154), .QN(n155) );
  NAND2X1 U330 ( .IN1(n614), .IN2(n527), .QN(n180) );
  NAND2X1 U331 ( .IN1(a_in[23]), .IN2(n316), .QN(n181) );
  NAND2X1 U332 ( .IN1(n609), .IN2(n463), .QN(n217) );
  NAND2X4 U333 ( .IN1(n302), .IN2(n312), .QN(n156) );
  NAND2X0 U334 ( .IN1(n541), .IN2(n540), .QN(n542) );
  INVX4 U335 ( .IN(n206), .QN(n160) );
  INVX8 U336 ( .IN(n160), .QN(n161) );
  NAND2X0 U337 ( .IN1(n614), .IN2(n465), .QN(n162) );
  NAND2X0 U338 ( .IN1(a_in[8]), .IN2(n319), .QN(n163) );
  NAND3X0 U339 ( .IN1(n162), .IN2(n163), .IN3(n129), .QN(N67) );
  NAND2X0 U340 ( .IN1(n614), .IN2(n583), .QN(n164) );
  NAND2X0 U341 ( .IN1(a_in[5]), .IN2(n314), .QN(n165) );
  NAND3X0 U342 ( .IN1(n164), .IN2(n165), .IN3(n130), .QN(N64) );
  NAND2X0 U343 ( .IN1(n614), .IN2(n561), .QN(n166) );
  NAND2X0 U344 ( .IN1(a_in[29]), .IN2(n315), .QN(n167) );
  NAND3X0 U345 ( .IN1(n166), .IN2(n167), .IN3(n121), .QN(N88) );
  NAND2X0 U346 ( .IN1(n614), .IN2(n567), .QN(n168) );
  NAND2X0 U347 ( .IN1(a_in[30]), .IN2(n315), .QN(n169) );
  NAND3X0 U348 ( .IN1(n168), .IN2(n169), .IN3(n122), .QN(N89) );
  NBUFFX16 U349 ( .IN(n612), .Q(n315) );
  NAND2X0 U350 ( .IN1(n614), .IN2(n468), .QN(n170) );
  NAND2X0 U351 ( .IN1(a_in[9]), .IN2(n319), .QN(n171) );
  NAND3X0 U352 ( .IN1(n170), .IN2(n171), .IN3(n123), .QN(N68) );
  NAND2X0 U353 ( .IN1(n614), .IN2(n613), .QN(n172) );
  NAND2X0 U354 ( .IN1(a_in[0]), .IN2(n313), .QN(n173) );
  NAND3X0 U355 ( .IN1(n172), .IN2(n173), .IN3(n131), .QN(N59) );
  NAND2X0 U356 ( .IN1(n614), .IN2(n518), .QN(n174) );
  NAND2X0 U357 ( .IN1(a_in[21]), .IN2(n316), .QN(n175) );
  NAND3X0 U358 ( .IN1(n174), .IN2(n175), .IN3(n128), .QN(N80) );
  NAND2X0 U359 ( .IN1(n614), .IN2(n530), .QN(n176) );
  NAND2X0 U360 ( .IN1(a_in[24]), .IN2(n313), .QN(n177) );
  NAND3X0 U361 ( .IN1(n176), .IN2(n177), .IN3(n125), .QN(N83) );
  NAND2X0 U362 ( .IN1(n614), .IN2(n491), .QN(n178) );
  NAND2X0 U363 ( .IN1(a_in[14]), .IN2(n317), .QN(n179) );
  NAND3X0 U364 ( .IN1(n178), .IN2(n179), .IN3(n124), .QN(N73) );
  NOR2X0 U365 ( .IN1(n423), .IN2(n422), .QN(n182) );
  NAND2X4 U366 ( .IN1(n186), .IN2(n185), .QN(n448) );
  OR2X1 U367 ( .IN1(n556), .IN2(n446), .Q(n185) );
  NOR2X4 U368 ( .IN1(n447), .IN2(n110), .QN(n186) );
  NAND2X2 U369 ( .IN1(n434), .IN2(n108), .QN(n435) );
  NAND3X0 U370 ( .IN1(n433), .IN2(n187), .IN3(n532), .QN(n539) );
  OR2X1 U371 ( .IN1(reg_b[27]), .IN2(n442), .Q(n190) );
  INVX1 U372 ( .IN(n287), .QN(n295) );
  OR4X1 U373 ( .IN1(n295), .IN2(n203), .IN3(reg_b[8]), .IN4(reg_b[9]), .Q(n59)
         );
  NAND2X4 U374 ( .IN1(n409), .IN2(n572), .QN(n411) );
  INVX16 U375 ( .IN(n600), .QN(n614) );
  INVX2 U376 ( .IN(n215), .QN(n288) );
  INVX0 U377 ( .IN(n194), .QN(n195) );
  NAND2X4 U378 ( .IN1(n207), .IN2(n208), .QN(n584) );
  NAND2X2 U379 ( .IN1(n569), .IN2(n573), .QN(n405) );
  AND2X2 U380 ( .IN1(n289), .IN2(n290), .Q(n228) );
  INVX2 U381 ( .IN(n260), .QN(n198) );
  INVX1 U382 ( .IN(n200), .QN(n201) );
  IBUFFX16 U383 ( .IN(n587), .QN(n589) );
  OR2X2 U384 ( .IN1(n295), .IN2(n413), .Q(n588) );
  NAND2X4 U385 ( .IN1(n411), .IN2(n410), .QN(n457) );
  NAND2X4 U386 ( .IN1(n453), .IN2(n115), .QN(n463) );
  OR2X2 U387 ( .IN1(n201), .IN2(n202), .Q(n419) );
  INVX2 U388 ( .IN(n460), .QN(n420) );
  NAND2X4 U389 ( .IN1(n418), .IN2(n417), .QN(n423) );
  NAND2X4 U390 ( .IN1(n250), .IN2(n112), .QN(n433) );
  INVX0 U391 ( .IN(n454), .QN(n456) );
  NOR2X0 U392 ( .IN1(n6), .IN2(n455), .QN(n259) );
  NAND2X0 U393 ( .IN1(n284), .IN2(n292), .QN(n208) );
  INVX4 U394 ( .IN(n580), .QN(n415) );
  INVX2 U395 ( .IN(n568), .QN(n406) );
  NAND2X4 U396 ( .IN1(n213), .IN2(n454), .QN(n609) );
  INVX0 U397 ( .IN(n455), .QN(n212) );
  AND2X2 U398 ( .IN1(n214), .IN2(n218), .Q(n219) );
  NAND2X4 U399 ( .IN1(n219), .IN2(n457), .QN(n418) );
  NAND2X4 U400 ( .IN1(n301), .IN2(n113), .QN(n250) );
  NAND2X4 U401 ( .IN1(n188), .IN2(n464), .QN(n600) );
  INVX0 U402 ( .IN(n517), .QN(n300) );
  NAND2X0 U403 ( .IN1(n279), .IN2(reg_a[21]), .QN(n520) );
  NOR2X4 U404 ( .IN1(n464), .IN2(n188), .QN(n220) );
  NOR2X4 U405 ( .IN1(n464), .IN2(n188), .QN(n221) );
  NOR2X4 U406 ( .IN1(n252), .IN2(n118), .QN(n226) );
  NOR2X4 U407 ( .IN1(n227), .IN2(n114), .QN(n252) );
  NOR2X4 U408 ( .IN1(n226), .IN2(n116), .QN(n225) );
  INVX0 U409 ( .IN(n400), .QN(n426) );
  NAND2X1 U410 ( .IN1(n261), .IN2(n204), .QN(n460) );
  OR2X1 U411 ( .IN1(reg_a[23]), .IN2(n389), .Q(n391) );
  NOR2X0 U412 ( .IN1(n541), .IN2(n111), .QN(n438) );
  NOR2X4 U413 ( .IN1(n423), .IN2(n422), .QN(n476) );
  INVX8 U414 ( .IN(n463), .QN(n464) );
  OA21X1 U415 ( .IN1(n533), .IN2(n255), .IN3(n532), .Q(n534) );
  OA21X1 U416 ( .IN1(n305), .IN2(n525), .IN3(n524), .Q(n526) );
  NAND2X0 U417 ( .IN1(n280), .IN2(reg_a[9]), .QN(n470) );
  NAND2X0 U418 ( .IN1(n273), .IN2(reg_b[21]), .QN(n519) );
  OAI21X1 U419 ( .IN1(reg_a[22]), .IN2(n281), .IN3(n519), .QN(n525) );
  NOR2X4 U420 ( .IN1(n251), .IN2(n117), .QN(n227) );
  NOR2X4 U421 ( .IN1(n464), .IN2(n188), .QN(n223) );
  NOR2X4 U422 ( .IN1(n464), .IN2(n188), .QN(n224) );
  NAND2X1 U423 ( .IN1(n550), .IN2(n549), .QN(N85) );
  NOR2X1 U424 ( .IN1(n548), .IN2(n547), .QN(n549) );
  OR3X2 U425 ( .IN1(n225), .IN2(n505), .IN3(n429), .Q(n430) );
  INVX0 U426 ( .IN(n525), .QN(n249) );
  NOR2X0 U427 ( .IN1(n308), .IN2(n517), .QN(n229) );
  AND2X1 U428 ( .IN1(n239), .IN2(n102), .Q(n407) );
  NAND2X0 U429 ( .IN1(reg_b[31]), .IN2(n230), .QN(n451) );
  XOR3X1 U430 ( .IN1(n277), .IN2(reg_a[10]), .IN3(n231), .Q(n473) );
  OAI21X1 U431 ( .IN1(n471), .IN2(n254), .IN3(n470), .QN(n231) );
  XOR3X1 U432 ( .IN1(n232), .IN2(reg_a[16]), .IN3(n233), .Q(n499) );
  OAI21X1 U433 ( .IN1(n497), .IN2(n258), .IN3(n496), .QN(n233) );
  XOR3X1 U434 ( .IN1(reg_b[19]), .IN2(n234), .IN3(n235), .Q(n512) );
  OAI21X1 U435 ( .IN1(n510), .IN2(n256), .IN3(n509), .QN(n235) );
  XOR3X1 U436 ( .IN1(reg_b[20]), .IN2(n236), .IN3(n237), .Q(n516) );
  OAI21X1 U437 ( .IN1(n515), .IN2(n514), .IN3(n513), .QN(n237) );
  XOR3X1 U438 ( .IN1(n281), .IN2(reg_a[22]), .IN3(n238), .Q(n523) );
  OAI21X1 U439 ( .IN1(n521), .IN2(n229), .IN3(n520), .QN(n238) );
  OR2X1 U440 ( .IN1(n239), .IN2(n102), .Q(n410) );
  OR2X1 U441 ( .IN1(reg_b[13]), .IN2(n240), .Q(n488) );
  OR2X1 U442 ( .IN1(reg_b[16]), .IN2(n241), .Q(n500) );
  NAND2X0 U443 ( .IN1(reg_b[28]), .IN2(n263), .QN(n443) );
  NOR2X4 U444 ( .IN1(n476), .IN2(n132), .QN(n251) );
  NBUFFX2 U445 ( .IN(n612), .Q(n319) );
  INVX0 U446 ( .IN(n345), .QN(n335) );
  INVX0 U447 ( .IN(n344), .QN(n337) );
  INVX0 U448 ( .IN(n345), .QN(n336) );
  INVX0 U449 ( .IN(n344), .QN(n338) );
  INVX0 U450 ( .IN(n312), .QN(n309) );
  INVX0 U451 ( .IN(n343), .QN(n340) );
  INVX0 U452 ( .IN(n342), .QN(n341) );
  INVX0 U453 ( .IN(n343), .QN(n339) );
  INVX0 U454 ( .IN(n321), .QN(n345) );
  INVX0 U455 ( .IN(n321), .QN(n344) );
  INVX0 U456 ( .IN(n6), .QN(n346) );
  INVX0 U457 ( .IN(n328), .QN(n347) );
  INVX0 U458 ( .IN(n322), .QN(n348) );
  INVX0 U459 ( .IN(n323), .QN(n350) );
  INVX0 U460 ( .IN(n323), .QN(n351) );
  INVX0 U461 ( .IN(n324), .QN(n352) );
  INVX0 U462 ( .IN(n324), .QN(n353) );
  INVX0 U463 ( .IN(n325), .QN(n354) );
  INVX0 U464 ( .IN(n325), .QN(n355) );
  INVX0 U465 ( .IN(n326), .QN(n356) );
  INVX0 U466 ( .IN(n326), .QN(n357) );
  INVX0 U467 ( .IN(n327), .QN(n358) );
  INVX0 U468 ( .IN(n322), .QN(n349) );
  INVX0 U469 ( .IN(n328), .QN(n361) );
  INVX0 U470 ( .IN(n327), .QN(n359) );
  INVX0 U471 ( .IN(n328), .QN(n360) );
  NOR2X0 U472 ( .IN1(n246), .IN2(n459), .QN(n244) );
  INVX0 U473 ( .IN(n588), .QN(n416) );
  INVX0 U474 ( .IN(n320), .QN(n342) );
  INVX0 U475 ( .IN(n333), .QN(n321) );
  INVX0 U476 ( .IN(n332), .QN(n322) );
  INVX0 U477 ( .IN(n332), .QN(n323) );
  INVX0 U478 ( .IN(n320), .QN(n343) );
  INVX0 U479 ( .IN(n331), .QN(n324) );
  INVX0 U480 ( .IN(n331), .QN(n325) );
  INVX0 U481 ( .IN(n330), .QN(n326) );
  INVX0 U482 ( .IN(n330), .QN(n327) );
  INVX0 U483 ( .IN(n329), .QN(n328) );
  OR2X1 U484 ( .IN1(n562), .IN2(n557), .Q(n446) );
  NOR2X0 U485 ( .IN1(n581), .IN2(n458), .QN(n246) );
  NOR2X0 U486 ( .IN1(n246), .IN2(n584), .QN(n247) );
  OR2X1 U487 ( .IN1(n557), .IN2(n564), .Q(n560) );
  OR2X1 U488 ( .IN1(n562), .IN2(n110), .Q(n566) );
  INVX0 U489 ( .IN(n509), .QN(n429) );
  NOR2X0 U490 ( .IN1(n603), .IN2(n602), .QN(n607) );
  NOR2X0 U491 ( .IN1(n599), .IN2(n598), .QN(n603) );
  NAND2X4 U492 ( .IN1(n134), .IN2(n294), .QN(n580) );
  INVX0 U493 ( .IN(n496), .QN(n427) );
  INVX0 U494 ( .IN(n484), .QN(n425) );
  NOR2X0 U495 ( .IN1(n545), .IN2(n544), .QN(n550) );
  NOR2X0 U496 ( .IN1(n599), .IN2(n536), .QN(n545) );
  INVX0 U497 ( .IN(n520), .QN(n432) );
  INVX0 U498 ( .IN(n6), .QN(n333) );
  INVX0 U499 ( .IN(n6), .QN(n332) );
  INVX0 U500 ( .IN(n6), .QN(n331) );
  INVX0 U501 ( .IN(n6), .QN(n330) );
  INVX0 U502 ( .IN(n6), .QN(n329) );
  INVX0 U503 ( .IN(n334), .QN(n320) );
  INVX0 U504 ( .IN(n6), .QN(n334) );
  INVX0 U505 ( .IN(n457), .QN(n581) );
  OR3X1 U506 ( .IN1(n283), .IN2(n616), .IN3(n615), .Q(gcd_ns[0]) );
  AND2X1 U507 ( .IN1(n212), .IN2(n326), .Q(n616) );
  OA21X1 U508 ( .IN1(n244), .IN2(n467), .IN3(n421), .Q(n254) );
  INVX0 U509 ( .IN(n537), .QN(n538) );
  INVX0 U510 ( .IN(n556), .QN(n564) );
  INVX0 U511 ( .IN(n563), .QN(n557) );
  INVX0 U512 ( .IN(n593), .QN(n562) );
  NOR2X0 U513 ( .IN1(n529), .IN2(n528), .QN(n255) );
  NOR2X0 U514 ( .IN1(n138), .IN2(n505), .QN(n256) );
  NOR2X0 U515 ( .IN1(n184), .IN2(n480), .QN(n257) );
  NOR2X0 U516 ( .IN1(n222), .IN2(n492), .QN(n258) );
  INVX0 U517 ( .IN(n394), .QN(n431) );
  INVX0 U518 ( .IN(n572), .QN(n574) );
  INVX0 U519 ( .IN(n469), .QN(n471) );
  INVX0 U520 ( .IN(n495), .QN(n497) );
  INVX0 U521 ( .IN(n508), .QN(n510) );
  INVX0 U522 ( .IN(n519), .QN(n521) );
  INVX0 U523 ( .IN(n531), .QN(n533) );
  INVX0 U524 ( .IN(n483), .QN(n485) );
  NBUFFX2 U525 ( .IN(n380), .Q(n375) );
  NBUFFX2 U526 ( .IN(n379), .Q(n377) );
  NBUFFX2 U527 ( .IN(n381), .Q(n374) );
  NBUFFX2 U528 ( .IN(n386), .Q(n363) );
  NBUFFX2 U529 ( .IN(n386), .Q(n364) );
  NBUFFX2 U530 ( .IN(n385), .Q(n365) );
  NBUFFX2 U531 ( .IN(n385), .Q(n366) );
  NBUFFX2 U532 ( .IN(n384), .Q(n367) );
  NBUFFX2 U533 ( .IN(n384), .Q(n368) );
  NBUFFX2 U534 ( .IN(n383), .Q(n369) );
  NBUFFX2 U535 ( .IN(n383), .Q(n370) );
  NBUFFX2 U536 ( .IN(n382), .Q(n371) );
  NBUFFX2 U537 ( .IN(n382), .Q(n372) );
  NBUFFX2 U538 ( .IN(n381), .Q(n373) );
  NBUFFX2 U539 ( .IN(n380), .Q(n376) );
  NBUFFX2 U540 ( .IN(n379), .Q(n378) );
  AO222X1 U541 ( .IN1(n615), .IN2(reg_a[31]), .IN3(b_in[31]), .IN4(n137), 
        .IN5(reg_b[31]), .IN6(n106), .Q(N123) );
  AO222X1 U542 ( .IN1(n103), .IN2(reg_a[20]), .IN3(b_in[20]), .IN4(n137), 
        .IN5(reg_b[20]), .IN6(n107), .Q(N112) );
  AO222X1 U543 ( .IN1(n104), .IN2(reg_a[22]), .IN3(b_in[22]), .IN4(n136), 
        .IN5(reg_b[22]), .IN6(n309), .Q(N114) );
  AO222X1 U544 ( .IN1(n103), .IN2(reg_a[23]), .IN3(b_in[23]), .IN4(n136), 
        .IN5(reg_b[23]), .IN6(n106), .Q(N115) );
  AO222X1 U545 ( .IN1(n615), .IN2(reg_a[10]), .IN3(b_in[10]), .IN4(n137), 
        .IN5(reg_b[10]), .IN6(n106), .Q(N102) );
  AO222X1 U546 ( .IN1(n103), .IN2(n195), .IN3(b_in[11]), .IN4(n136), .IN5(
        reg_b[11]), .IN6(n107), .Q(N103) );
  AO222X1 U547 ( .IN1(n615), .IN2(reg_a[14]), .IN3(b_in[14]), .IN4(n137), 
        .IN5(reg_b[14]), .IN6(n107), .Q(N106) );
  AO222X1 U548 ( .IN1(n103), .IN2(reg_a[15]), .IN3(b_in[15]), .IN4(n137), 
        .IN5(reg_b[15]), .IN6(n107), .Q(N107) );
  AO222X1 U549 ( .IN1(n303), .IN2(reg_a[16]), .IN3(b_in[16]), .IN4(n137), 
        .IN5(reg_b[16]), .IN6(n309), .Q(N108) );
  AO222X1 U550 ( .IN1(n303), .IN2(reg_a[17]), .IN3(b_in[17]), .IN4(n136), 
        .IN5(reg_b[17]), .IN6(n106), .Q(N109) );
  AO222X1 U551 ( .IN1(n104), .IN2(reg_a[25]), .IN3(b_in[25]), .IN4(n137), 
        .IN5(reg_b[25]), .IN6(n107), .Q(N117) );
  AO222X1 U552 ( .IN1(n103), .IN2(reg_a[27]), .IN3(b_in[27]), .IN4(n137), 
        .IN5(reg_b[27]), .IN6(n106), .Q(N119) );
  AO222X1 U553 ( .IN1(n615), .IN2(reg_a[29]), .IN3(b_in[29]), .IN4(n136), 
        .IN5(reg_b[29]), .IN6(n106), .Q(N121) );
  AO222X1 U554 ( .IN1(n615), .IN2(reg_a[3]), .IN3(b_in[3]), .IN4(n137), .IN5(
        n102), .IN6(n107), .Q(N95) );
  NAND2X0 U555 ( .IN1(n260), .IN2(reg_b[2]), .QN(n572) );
  AND3X1 U556 ( .IN1(reg_a[31]), .IN2(n595), .IN3(n594), .Q(n597) );
  OAI21X1 U557 ( .IN1(n110), .IN2(n248), .IN3(n593), .QN(n594) );
  MUX21X1 U558 ( .IN1(n560), .IN2(n559), .S(n148), .Q(n561) );
  XOR2X1 U559 ( .IN1(n274), .IN2(reg_a[29]), .Q(n559) );
  XOR3X1 U560 ( .IN1(n102), .IN2(reg_a[3]), .IN3(n575), .Q(n577) );
  OA21X1 U561 ( .IN1(n574), .IN2(n253), .IN3(n573), .Q(n575) );
  XOR3X1 U562 ( .IN1(reg_b[25]), .IN2(reg_a[25]), .IN3(n534), .Q(n535) );
  XOR3X1 U563 ( .IN1(reg_a[2]), .IN2(reg_b[2]), .IN3(n253), .Q(n571) );
  XOR3X1 U564 ( .IN1(reg_b[23]), .IN2(reg_a[23]), .IN3(n526), .Q(n527) );
  AND2X1 U565 ( .IN1(reg_b[1]), .IN2(n221), .Q(n604) );
  AND2X1 U566 ( .IN1(reg_b[26]), .IN2(n220), .Q(n547) );
  MUX21X1 U567 ( .IN1(n566), .IN2(n565), .S(n248), .Q(n567) );
  XOR2X1 U568 ( .IN1(n275), .IN2(reg_a[30]), .Q(n565) );
  XOR3X1 U569 ( .IN1(reg_a[12]), .IN2(reg_b[12]), .IN3(n257), .Q(n482) );
  XOR3X1 U570 ( .IN1(reg_a[15]), .IN2(reg_b[15]), .IN3(n258), .Q(n494) );
  XOR3X1 U571 ( .IN1(reg_a[18]), .IN2(reg_b[18]), .IN3(n256), .Q(n507) );
  XOR3X1 U572 ( .IN1(reg_a[21]), .IN2(reg_b[21]), .IN3(n229), .Q(n518) );
  XOR3X1 U573 ( .IN1(reg_a[24]), .IN2(reg_b[24]), .IN3(n255), .Q(n530) );
  OA21X1 U574 ( .IN1(n485), .IN2(n257), .IN3(n484), .Q(n486) );
  OA21X1 U575 ( .IN1(n589), .IN2(n247), .IN3(n588), .Q(n590) );
  XOR3X1 U576 ( .IN1(reg_b[17]), .IN2(reg_a[17]), .IN3(n502), .Q(n504) );
  OAI21X1 U577 ( .IN1(reg_b[0]), .IN2(n611), .IN3(n610), .QN(n613) );
  INVX0 U578 ( .IN(reg_a[0]), .QN(n611) );
  XOR3X1 U579 ( .IN1(reg_b[26]), .IN2(reg_a[26]), .IN3(n542), .Q(n543) );
  XOR3X1 U580 ( .IN1(n296), .IN2(n610), .IN3(reg_b[1]), .Q(n601) );
  OAI21X1 U581 ( .IN1(reg_a[25]), .IN2(n278), .IN3(n531), .QN(n537) );
  AO22X1 U582 ( .IN1(n390), .IN2(n391), .IN3(reg_a[23]), .IN4(n389), .Q(n528)
         );
  AO22X1 U583 ( .IN1(n399), .IN2(n400), .IN3(reg_a[14]), .IN4(n398), .Q(n492)
         );
  INVX0 U584 ( .IN(n488), .QN(n399) );
  AO22X1 U585 ( .IN1(n402), .IN2(n403), .IN3(reg_a[11]), .IN4(n191), .Q(n480)
         );
  INVX0 U586 ( .IN(n474), .QN(n402) );
  OR4X1 U587 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n63) );
  OR4X1 U588 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n62) );
  OR4X1 U589 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(
        reg_b[16]), .Q(n65) );
  OR2X1 U590 ( .IN1(reg_a[29]), .IN2(n274), .Q(n556) );
  AO22X1 U591 ( .IN1(reg_a[8]), .IN2(n346), .IN3(result[8]), .IN4(n322), .Q(
        n68) );
  AO22X1 U592 ( .IN1(reg_a[9]), .IN2(n347), .IN3(result[9]), .IN4(n341), .Q(
        n69) );
  AO22X1 U593 ( .IN1(reg_a[10]), .IN2(n347), .IN3(result[10]), .IN4(n341), .Q(
        n70) );
  AO22X1 U594 ( .IN1(n195), .IN2(n348), .IN3(result[11]), .IN4(n341), .Q(n71)
         );
  AO22X1 U595 ( .IN1(reg_a[12]), .IN2(n348), .IN3(result[12]), .IN4(n341), .Q(
        n72) );
  AO22X1 U596 ( .IN1(reg_a[14]), .IN2(n349), .IN3(result[14]), .IN4(n340), .Q(
        n74) );
  AO22X1 U597 ( .IN1(reg_a[15]), .IN2(n350), .IN3(result[15]), .IN4(n340), .Q(
        n75) );
  AO22X1 U598 ( .IN1(reg_a[16]), .IN2(n350), .IN3(result[16]), .IN4(n340), .Q(
        n76) );
  AO22X1 U599 ( .IN1(reg_a[17]), .IN2(n351), .IN3(result[17]), .IN4(n339), .Q(
        n77) );
  AO22X1 U600 ( .IN1(reg_a[18]), .IN2(n351), .IN3(result[18]), .IN4(n339), .Q(
        n78) );
  AO22X1 U601 ( .IN1(reg_a[19]), .IN2(n352), .IN3(result[19]), .IN4(n339), .Q(
        n79) );
  AO22X1 U602 ( .IN1(reg_a[20]), .IN2(n352), .IN3(result[20]), .IN4(n339), .Q(
        n80) );
  AO22X1 U603 ( .IN1(reg_a[21]), .IN2(n353), .IN3(result[21]), .IN4(n338), .Q(
        n81) );
  AO22X1 U604 ( .IN1(reg_a[22]), .IN2(n353), .IN3(result[22]), .IN4(n338), .Q(
        n82) );
  AO22X1 U605 ( .IN1(reg_a[23]), .IN2(n354), .IN3(result[23]), .IN4(n338), .Q(
        n83) );
  AO22X1 U606 ( .IN1(reg_a[24]), .IN2(n354), .IN3(result[24]), .IN4(n337), .Q(
        n84) );
  AO22X1 U607 ( .IN1(reg_a[25]), .IN2(n355), .IN3(result[25]), .IN4(n337), .Q(
        n85) );
  AO22X1 U608 ( .IN1(reg_a[26]), .IN2(n355), .IN3(result[26]), .IN4(n337), .Q(
        n86) );
  AO22X1 U609 ( .IN1(reg_a[27]), .IN2(n356), .IN3(result[27]), .IN4(n337), .Q(
        n87) );
  AO22X1 U610 ( .IN1(reg_a[28]), .IN2(n356), .IN3(result[28]), .IN4(n336), .Q(
        n88) );
  AO22X1 U611 ( .IN1(reg_a[29]), .IN2(n357), .IN3(result[29]), .IN4(n336), .Q(
        n89) );
  AO22X1 U612 ( .IN1(reg_a[30]), .IN2(n357), .IN3(result[30]), .IN4(n336), .Q(
        n90) );
  AO22X1 U613 ( .IN1(reg_a[2]), .IN2(n358), .IN3(result[2]), .IN4(n336), .Q(
        n91) );
  AO22X1 U614 ( .IN1(reg_a[3]), .IN2(n358), .IN3(result[3]), .IN4(n335), .Q(
        n92) );
  AO22X1 U615 ( .IN1(reg_a[31]), .IN2(n361), .IN3(result[31]), .IN4(n327), .Q(
        n97) );
  AO22X1 U616 ( .IN1(reg_a[0]), .IN2(n347), .IN3(result[0]), .IN4(n338), .Q(
        n99) );
  OR2X2 U617 ( .IN1(reg_a[11]), .IN2(n191), .Q(n403) );
  NAND2X0 U618 ( .IN1(n269), .IN2(reg_a[24]), .QN(n532) );
  NAND2X0 U619 ( .IN1(n274), .IN2(reg_a[29]), .QN(n563) );
  NAND2X0 U620 ( .IN1(n275), .IN2(reg_a[30]), .QN(n593) );
  NAND2X0 U621 ( .IN1(reg_a[26]), .IN2(n388), .QN(n436) );
  NAND2X0 U622 ( .IN1(reg_a[31]), .IN2(n595), .QN(n449) );
  NAND2X0 U623 ( .IN1(n278), .IN2(reg_a[25]), .QN(n541) );
  NAND2X0 U624 ( .IN1(reg_b[27]), .IN2(n442), .QN(n440) );
  OAI21X1 U625 ( .IN1(reg_a[16]), .IN2(n232), .IN3(n495), .QN(n501) );
  INVX0 U626 ( .IN(a_in[1]), .QN(n598) );
  INVX0 U627 ( .IN(a_in[26]), .QN(n536) );
  NAND2X0 U628 ( .IN1(n281), .IN2(reg_a[22]), .QN(n524) );
  AND2X1 U629 ( .IN1(n282), .IN2(n67), .Q(done) );
  AND3X1 U630 ( .IN1(start), .IN2(n67), .IN3(n100), .Q(n283) );
  AO22X1 U631 ( .IN1(n396), .IN2(n397), .IN3(reg_a[17]), .IN4(n395), .Q(n505)
         );
  NBUFFX2 U632 ( .IN(n387), .Q(n362) );
  NBUFFX2 U633 ( .IN(reset_n), .Q(n387) );
  NBUFFX2 U634 ( .IN(reset_n), .Q(n386) );
  NBUFFX2 U635 ( .IN(reset_n), .Q(n385) );
  NBUFFX2 U636 ( .IN(reset_n), .Q(n384) );
  NBUFFX2 U637 ( .IN(reset_n), .Q(n383) );
  NBUFFX2 U638 ( .IN(reset_n), .Q(n382) );
  NBUFFX2 U639 ( .IN(reset_n), .Q(n381) );
  NBUFFX2 U640 ( .IN(reset_n), .Q(n380) );
  NBUFFX2 U641 ( .IN(reset_n), .Q(n379) );
  XOR3X1 U642 ( .IN1(reg_b[13]), .IN2(reg_a[13]), .IN3(n486), .Q(n487) );
  OAI21X1 U643 ( .IN1(reg_a[13]), .IN2(n401), .IN3(n483), .QN(n489) );
  AO22X1 U644 ( .IN1(reg_a[13]), .IN2(n349), .IN3(result[13]), .IN4(n340), .Q(
        n73) );
  AO222X1 U645 ( .IN1(n104), .IN2(n204), .IN3(b_in[7]), .IN4(n136), .IN5(n203), 
        .IN6(n309), .Q(N99) );
  AO22X1 U646 ( .IN1(n204), .IN2(n360), .IN3(result[7]), .IN4(n324), .Q(n96)
         );
  INVX0 U647 ( .IN(n312), .QN(n311) );
  AO22X1 U648 ( .IN1(n296), .IN2(n361), .IN3(result[1]), .IN4(n325), .Q(n98)
         );
  OA21X1 U649 ( .IN1(n244), .IN2(n461), .IN3(n460), .Q(n462) );
  OA21X1 U650 ( .IN1(n581), .IN2(n228), .IN3(n580), .Q(n582) );
  NOR2X0 U651 ( .IN1(n601), .IN2(n600), .QN(n602) );
  NOR2X0 U652 ( .IN1(n543), .IN2(n600), .QN(n544) );
  AO222X1 U653 ( .IN1(n103), .IN2(reg_a[2]), .IN3(b_in[2]), .IN4(n136), .IN5(
        reg_b[2]), .IN6(n106), .Q(N94) );
  OR4X1 U654 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n61) );
  AO221X1 U655 ( .IN1(n614), .IN2(n523), .IN3(a_in[22]), .IN4(n319), .IN5(n522), .Q(N81) );
  AO222X1 U656 ( .IN1(n303), .IN2(reg_a[30]), .IN3(b_in[30]), .IN4(n137), 
        .IN5(reg_b[30]), .IN6(n107), .Q(N122) );
  AO222X1 U657 ( .IN1(n103), .IN2(reg_a[24]), .IN3(b_in[24]), .IN4(n137), 
        .IN5(reg_b[24]), .IN6(n311), .Q(N116) );
  AO222X1 U658 ( .IN1(n104), .IN2(reg_a[19]), .IN3(b_in[19]), .IN4(n137), 
        .IN5(reg_b[19]), .IN6(n309), .Q(N111) );
  AO222X1 U659 ( .IN1(n615), .IN2(reg_a[12]), .IN3(b_in[12]), .IN4(n137), 
        .IN5(reg_b[12]), .IN6(n106), .Q(N104) );
  INVX8 U660 ( .IN(n609), .QN(n312) );
  AO22X1 U661 ( .IN1(n420), .IN2(n419), .IN3(reg_a[8]), .IN4(n202), .Q(n466)
         );
  OR4X1 U662 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(
        reg_b[1]), .Q(n64) );
  NAND2X0 U663 ( .IN1(n539), .IN2(n538), .QN(n540) );
  AO22X1 U664 ( .IN1(n284), .IN2(n359), .IN3(result[5]), .IN4(n335), .Q(n94)
         );
  AO22X1 U665 ( .IN1(n288), .IN2(n360), .IN3(result[6]), .IN4(n335), .Q(n95)
         );
  OR4X1 U666 ( .IN1(reg_b[31]), .IN2(n102), .IN3(n290), .IN4(n293), .Q(n60) );
  AO222X1 U667 ( .IN1(n615), .IN2(n294), .IN3(b_in[4]), .IN4(n136), .IN5(n290), 
        .IN6(n107), .Q(N96) );
  XOR3X1 U668 ( .IN1(n294), .IN2(n290), .IN3(n581), .Q(n579) );
  AO22X1 U669 ( .IN1(n294), .IN2(n359), .IN3(result[4]), .IN4(n335), .Q(n93)
         );
  INVX2 U670 ( .IN(n298), .QN(n299) );
  AO221X1 U671 ( .IN1(n614), .IN2(n504), .IN3(a_in[17]), .IN4(n317), .IN5(n503), .Q(N76) );
  AO222X1 U672 ( .IN1(n303), .IN2(reg_a[9]), .IN3(b_in[9]), .IN4(n136), .IN5(
        reg_b[9]), .IN6(n107), .Q(N101) );
  AO222X1 U673 ( .IN1(n103), .IN2(reg_a[21]), .IN3(b_in[21]), .IN4(n136), 
        .IN5(reg_b[21]), .IN6(n106), .Q(N113) );
  AO222X1 U674 ( .IN1(n104), .IN2(reg_a[18]), .IN3(b_in[18]), .IN4(n136), 
        .IN5(reg_b[18]), .IN6(n311), .Q(N110) );
  AO222X1 U675 ( .IN1(n104), .IN2(reg_a[28]), .IN3(b_in[28]), .IN4(n136), 
        .IN5(reg_b[28]), .IN6(n311), .Q(N120) );
  AO222X1 U676 ( .IN1(n104), .IN2(n284), .IN3(b_in[5]), .IN4(n136), .IN5(n293), 
        .IN6(n311), .Q(N97) );
  AO222X1 U677 ( .IN1(n104), .IN2(n296), .IN3(b_in[1]), .IN4(n136), .IN5(
        reg_b[1]), .IN6(n106), .Q(N93) );
  AO222X1 U678 ( .IN1(n104), .IN2(reg_a[26]), .IN3(b_in[26]), .IN4(n136), 
        .IN5(reg_b[26]), .IN6(n106), .Q(N118) );
  AO222X1 U679 ( .IN1(n615), .IN2(reg_a[13]), .IN3(b_in[13]), .IN4(n136), 
        .IN5(reg_b[13]), .IN6(n309), .Q(N105) );
  AO222X1 U680 ( .IN1(n103), .IN2(reg_a[8]), .IN3(b_in[8]), .IN4(n137), .IN5(
        reg_b[8]), .IN6(n107), .Q(N100) );
  NOR2X0 U681 ( .IN1(n546), .IN2(n291), .QN(n548) );
  NAND2X4 U682 ( .IN1(n464), .IN2(n312), .QN(n599) );
  AND2X1 U683 ( .IN1(n259), .IN2(n159), .Q(gcd_ns[1]) );
  AND3X1 U684 ( .IN1(n394), .IN2(n306), .IN3(n430), .Q(n304) );
  NOR3X0 U685 ( .IN1(n304), .IN2(n517), .IN3(n432), .QN(n305) );
  NOR3X0 U686 ( .IN1(n431), .IN2(n514), .IN3(n515), .QN(n308) );
  AO221X1 U687 ( .IN1(n614), .IN2(n499), .IN3(a_in[16]), .IN4(n317), .IN5(n498), .Q(N75) );
  AO221X1 U688 ( .IN1(n614), .IN2(n555), .IN3(a_in[28]), .IN4(n315), .IN5(n554), .Q(N87) );
  AO221X1 U689 ( .IN1(n614), .IN2(n577), .IN3(a_in[3]), .IN4(n314), .IN5(n576), 
        .Q(N62) );
  AO22X1 U690 ( .IN1(n221), .IN2(reg_b[12]), .IN3(n285), .IN4(reg_a[12]), .Q(
        n481) );
  AO221X1 U691 ( .IN1(n614), .IN2(n479), .IN3(a_in[11]), .IN4(n318), .IN5(n478), .Q(N70) );
  AO22X1 U692 ( .IN1(n220), .IN2(reg_b[11]), .IN3(n161), .IN4(n195), .Q(n478)
         );
  AO221X1 U693 ( .IN1(n614), .IN2(n512), .IN3(a_in[19]), .IN4(n316), .IN5(n511), .Q(N78) );
  AO22X1 U694 ( .IN1(n220), .IN2(reg_b[19]), .IN3(n161), .IN4(reg_a[19]), .Q(
        n511) );
  AO221X1 U695 ( .IN1(n614), .IN2(n507), .IN3(a_in[18]), .IN4(n316), .IN5(n506), .Q(N77) );
  AO22X1 U696 ( .IN1(n221), .IN2(reg_b[18]), .IN3(n161), .IN4(reg_a[18]), .Q(
        n506) );
  AO221X1 U697 ( .IN1(n614), .IN2(n494), .IN3(a_in[15]), .IN4(n317), .IN5(n493), .Q(N74) );
  AO22X1 U698 ( .IN1(n223), .IN2(reg_b[15]), .IN3(n285), .IN4(reg_a[15]), .Q(
        n493) );
  AO221X1 U699 ( .IN1(n614), .IN2(n473), .IN3(a_in[10]), .IN4(n318), .IN5(n472), .Q(N69) );
  AO22X1 U700 ( .IN1(n223), .IN2(reg_b[10]), .IN3(n285), .IN4(reg_a[10]), .Q(
        n472) );
  AO22X1 U701 ( .IN1(n224), .IN2(n290), .IN3(n161), .IN4(n294), .Q(n578) );
  OA21X1 U702 ( .IN1(n139), .IN2(n501), .IN3(n500), .Q(n502) );
  AO221X1 U703 ( .IN1(n614), .IN2(n579), .IN3(a_in[4]), .IN4(n314), .IN5(n578), 
        .Q(N63) );
  AO22X1 U704 ( .IN1(n224), .IN2(reg_b[31]), .IN3(n161), .IN4(reg_a[31]), .Q(
        n596) );
  AO221X1 U705 ( .IN1(n614), .IN2(n553), .IN3(a_in[27]), .IN4(n315), .IN5(n552), .Q(N86) );
  AO22X1 U706 ( .IN1(n223), .IN2(reg_b[27]), .IN3(n285), .IN4(reg_a[27]), .Q(
        n552) );
  AO221X1 U707 ( .IN1(n614), .IN2(n592), .IN3(a_in[7]), .IN4(n313), .IN5(n591), 
        .Q(N66) );
  AO22X1 U708 ( .IN1(n224), .IN2(n203), .IN3(n161), .IN4(n204), .Q(n591) );
  AO221X1 U709 ( .IN1(n614), .IN2(n571), .IN3(a_in[2]), .IN4(n314), .IN5(n570), 
        .Q(N61) );
  AO22X1 U710 ( .IN1(n223), .IN2(reg_b[2]), .IN3(n161), .IN4(reg_a[2]), .Q(
        n570) );
  AO22X1 U711 ( .IN1(n223), .IN2(reg_b[16]), .IN3(n161), .IN4(reg_a[16]), .Q(
        n498) );
  AO22X1 U712 ( .IN1(n220), .IN2(reg_b[17]), .IN3(n285), .IN4(reg_a[17]), .Q(
        n503) );
  OA21X1 U713 ( .IN1(n183), .IN2(n489), .IN3(n488), .Q(n490) );
  AO222X1 U714 ( .IN1(reg_a[0]), .IN2(n303), .IN3(b_in[0]), .IN4(n137), .IN5(
        reg_b[0]), .IN6(n311), .Q(N92) );
  AO221X1 U715 ( .IN1(n614), .IN2(n586), .IN3(a_in[6]), .IN4(n313), .IN5(n585), 
        .Q(N65) );
  AO22X1 U716 ( .IN1(n224), .IN2(n295), .IN3(n285), .IN4(n288), .Q(n585) );
  AO22X1 U717 ( .IN1(n221), .IN2(reg_b[22]), .IN3(n161), .IN4(reg_a[22]), .Q(
        n522) );
  AO221X1 U718 ( .IN1(n614), .IN2(n482), .IN3(a_in[12]), .IN4(n318), .IN5(n481), .Q(N71) );
  OA21X1 U719 ( .IN1(n182), .IN2(n475), .IN3(n474), .Q(n477) );
  AO221X1 U720 ( .IN1(n614), .IN2(n597), .IN3(a_in[31]), .IN4(n313), .IN5(n596), .Q(N90) );
  AO22X1 U721 ( .IN1(n223), .IN2(reg_b[28]), .IN3(n285), .IN4(reg_a[28]), .Q(
        n554) );
  AO22X1 U722 ( .IN1(n224), .IN2(n102), .IN3(n285), .IN4(reg_a[3]), .Q(n576)
         );
  INVX4 U723 ( .IN(n551), .QN(n439) );
  OR2X2 U724 ( .IN1(n299), .IN2(n307), .Q(n610) );
  NAND2X4 U725 ( .IN1(n435), .IN2(n436), .QN(n437) );
  NOR2X4 U726 ( .IN1(n438), .IN2(n437), .QN(n551) );
  NAND2X4 U727 ( .IN1(n439), .IN2(n440), .QN(n441) );
  NAND2X4 U728 ( .IN1(n445), .IN2(n444), .QN(n558) );
  NOR2X4 U729 ( .IN1(n558), .IN2(n446), .QN(n447) );
  NAND2X4 U730 ( .IN1(n450), .IN2(n451), .QN(n452) );
  INVX8 U731 ( .IN(n599), .QN(n612) );
endmodule

