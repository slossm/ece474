library verilog;
use verilog.vl_types.all;
entity stoplighttb is
    generic(
        CYCLE           : integer := 100
    );
end stoplighttb;
